magic
tech scmos
timestamp 1085807705
<< polysilicon >>
rect 37 429 40 497
rect 45 855 3722 857
rect 45 850 3722 852
rect 45 845 3722 847
rect 45 840 3722 842
rect 45 835 3722 837
rect 45 830 3722 832
rect 45 825 3722 827
rect 45 820 3722 822
rect 45 815 3722 817
rect 45 810 3722 812
rect 45 805 3722 807
rect 45 800 3722 802
rect 45 795 3722 797
rect 45 790 3722 792
rect 45 785 3722 787
rect 45 780 3722 782
rect 45 775 3722 777
rect 45 770 3722 772
rect 45 765 3722 767
rect 45 760 3722 762
rect 45 755 3722 757
rect 45 750 3722 752
rect 45 745 3722 747
rect 45 740 3722 742
rect 45 735 3722 737
rect 45 730 3722 732
rect 45 725 3722 727
rect 45 720 3722 722
rect 45 715 3722 717
rect 45 710 3722 712
rect 45 705 3722 707
rect 45 700 3722 702
rect 45 695 3722 697
rect 45 690 3722 692
rect 45 685 3722 687
rect 45 680 3722 682
rect 45 675 3722 677
rect 45 670 3722 672
rect 45 665 3722 667
rect 45 660 3722 662
rect 45 655 3722 657
rect 45 650 3722 652
rect 45 645 3722 647
rect 45 640 3722 642
rect 45 635 3722 637
rect 45 630 3722 632
rect 45 625 3722 627
rect 45 620 3722 622
rect 45 615 3722 617
rect 45 610 3722 612
rect 45 605 3722 607
rect 45 600 3722 602
rect 45 595 3722 597
rect 45 590 3722 592
rect 45 585 3722 587
rect 45 580 3722 582
rect 45 575 3722 577
rect 45 570 3722 572
rect 45 565 3722 567
rect 45 560 3722 562
rect 45 555 3722 557
rect 45 550 3722 552
rect 45 545 3722 547
rect 45 540 3722 542
rect 45 535 3722 537
rect 45 530 3722 532
rect 45 525 3722 527
rect 45 520 3722 522
rect 45 515 3722 517
rect 45 510 3722 512
rect 45 505 3722 507
rect 45 500 3722 502
rect 45 495 3722 497
rect 45 490 3722 492
rect 45 485 3722 487
rect 45 480 3722 482
rect 45 475 3722 477
rect 45 470 3722 472
rect 45 465 3722 467
rect 45 460 3722 462
rect 45 455 3722 457
rect 45 450 3722 452
rect 45 445 3722 447
rect 45 440 3722 442
rect 45 435 3722 437
rect 45 430 3722 432
rect 45 425 3722 427
rect 45 420 3722 422
rect 45 415 3722 417
rect 45 410 3722 412
rect 45 405 3722 407
rect 45 400 3722 402
rect 45 395 3722 397
rect 45 390 3722 392
rect 45 385 3722 387
rect 45 380 3722 382
rect 45 375 3722 377
rect 45 370 3722 372
rect 45 365 3722 367
rect 45 360 3722 362
rect 45 355 3722 357
rect 45 350 3722 352
rect 45 345 3722 347
rect 45 340 3722 342
rect 45 335 3722 337
rect 45 330 3722 332
rect 45 325 3722 327
rect 45 320 3722 322
rect 45 315 3722 317
rect 45 310 3722 312
rect 45 305 3722 307
rect 45 300 3722 302
rect 45 295 3722 297
rect 45 290 3722 292
rect 45 285 3722 287
rect 45 280 3722 282
rect 45 275 3722 277
rect 45 270 3722 272
rect 45 265 3722 267
rect 45 260 3722 262
rect 45 255 3722 257
rect 45 250 3722 252
rect 45 245 3722 247
rect 45 240 3722 242
rect 45 235 3722 237
rect 45 230 3722 232
rect 45 225 3722 227
rect 45 220 3722 222
rect 45 215 3722 217
rect 45 210 3722 212
rect 45 205 3722 207
rect 45 200 3722 202
rect 45 195 3722 197
rect 45 190 3722 192
rect 45 185 3722 187
rect 45 180 3722 182
rect 45 175 3722 177
rect 45 170 3722 172
rect 45 165 3722 167
rect 45 160 3722 162
rect 45 155 3722 157
rect 45 150 3722 152
rect 45 145 3722 147
rect 45 140 3722 142
rect 45 135 3722 137
rect 45 130 3722 132
rect 45 125 3722 127
rect 45 120 3722 122
rect 45 115 3722 117
rect 45 110 3722 112
rect 45 105 3722 107
rect 45 100 3722 102
rect 45 95 3722 97
rect 45 90 3722 92
rect 45 85 3722 87
rect 45 80 3722 82
rect 45 75 3722 77
rect 45 70 3722 72
rect 45 65 3722 67
rect 45 60 3722 62
<< metal1 >>
rect 37 429 40 497
rect 45 855 60 857
rect 45 850 3722 855
rect 45 845 60 850
rect 45 840 3722 845
rect 45 835 60 840
rect 45 830 3722 835
rect 45 825 60 830
rect 45 820 3722 825
rect 45 815 60 820
rect 45 810 3722 815
rect 45 805 60 810
rect 45 800 3722 805
rect 45 795 60 800
rect 45 790 3722 795
rect 45 785 60 790
rect 45 780 3722 785
rect 45 775 60 780
rect 45 770 3722 775
rect 45 765 60 770
rect 45 760 3722 765
rect 45 755 60 760
rect 45 750 3722 755
rect 45 745 60 750
rect 45 740 3722 745
rect 45 735 60 740
rect 45 730 3722 735
rect 45 725 60 730
rect 45 720 3722 725
rect 45 715 60 720
rect 45 710 3722 715
rect 45 705 60 710
rect 45 700 3722 705
rect 45 695 60 700
rect 45 690 3722 695
rect 45 685 60 690
rect 45 680 3722 685
rect 45 675 60 680
rect 45 670 3722 675
rect 45 665 60 670
rect 45 660 3722 665
rect 45 655 60 660
rect 45 650 3722 655
rect 45 645 60 650
rect 45 640 3722 645
rect 45 635 60 640
rect 45 630 3722 635
rect 45 625 60 630
rect 45 620 3722 625
rect 45 615 60 620
rect 45 610 3722 615
rect 45 605 60 610
rect 45 600 3722 605
rect 45 595 60 600
rect 45 590 3722 595
rect 45 585 60 590
rect 45 580 3722 585
rect 45 575 60 580
rect 45 570 3722 575
rect 45 565 60 570
rect 45 560 3722 565
rect 45 555 60 560
rect 45 550 3722 555
rect 45 545 60 550
rect 45 540 3722 545
rect 45 535 60 540
rect 45 530 3722 535
rect 45 525 60 530
rect 45 520 3722 525
rect 45 515 60 520
rect 45 510 3722 515
rect 45 505 60 510
rect 45 500 3722 505
rect 45 495 60 500
rect 45 490 3722 495
rect 45 485 60 490
rect 45 480 3722 485
rect 45 475 60 480
rect 45 470 3722 475
rect 45 465 60 470
rect 45 460 3722 465
rect 45 455 60 460
rect 45 450 3722 455
rect 45 445 60 450
rect 45 440 3722 445
rect 45 435 60 440
rect 45 430 3722 435
rect 45 425 60 430
rect 45 420 3722 425
rect 45 415 60 420
rect 45 410 3722 415
rect 45 405 60 410
rect 45 400 3722 405
rect 45 395 60 400
rect 45 390 3722 395
rect 45 385 60 390
rect 45 380 3722 385
rect 45 375 60 380
rect 45 370 3722 375
rect 45 365 60 370
rect 45 360 3722 365
rect 45 355 60 360
rect 45 350 3722 355
rect 45 345 60 350
rect 45 340 3722 345
rect 45 335 60 340
rect 45 330 3722 335
rect 45 325 60 330
rect 45 320 3722 325
rect 45 315 60 320
rect 45 310 3722 315
rect 45 305 60 310
rect 45 300 3722 305
rect 45 295 60 300
rect 45 290 3722 295
rect 45 285 60 290
rect 45 280 3722 285
rect 45 275 60 280
rect 45 270 3722 275
rect 45 265 60 270
rect 45 260 3722 265
rect 45 255 60 260
rect 45 250 3722 255
rect 45 245 60 250
rect 45 240 3722 245
rect 45 235 60 240
rect 45 230 3722 235
rect 45 225 60 230
rect 45 220 3722 225
rect 45 215 60 220
rect 45 210 3722 215
rect 45 205 60 210
rect 45 200 3722 205
rect 45 195 60 200
rect 45 190 3722 195
rect 45 185 60 190
rect 45 180 3722 185
rect 45 175 60 180
rect 45 170 3722 175
rect 45 165 60 170
rect 45 160 3722 165
rect 45 155 60 160
rect 45 150 3722 155
rect 45 145 60 150
rect 45 140 3722 145
rect 45 135 60 140
rect 45 130 3722 135
rect 45 125 60 130
rect 45 120 3722 125
rect 45 115 60 120
rect 45 110 3722 115
rect 45 105 60 110
rect 45 100 3722 105
rect 45 95 60 100
rect 45 90 3722 95
rect 45 85 60 90
rect 45 80 3722 85
rect 45 75 60 80
rect 45 70 3722 75
rect 45 65 60 70
rect 45 60 3722 65
<< pm12contact >>
rect 29 429 37 497
rect 40 60 45 857
<< metal2 >>
rect 28 429 29 497
rect 37 429 40 497
rect 45 60 46 857
rect 51 855 60 857
rect 51 850 3722 855
rect 51 845 60 850
rect 51 840 3722 845
rect 51 835 60 840
rect 51 830 3722 835
rect 51 825 60 830
rect 51 820 3722 825
rect 51 815 60 820
rect 51 810 3722 815
rect 51 805 60 810
rect 51 800 3722 805
rect 51 795 60 800
rect 51 790 3722 795
rect 51 785 60 790
rect 51 780 3722 785
rect 51 775 60 780
rect 51 770 3722 775
rect 51 765 60 770
rect 51 760 3722 765
rect 51 755 60 760
rect 51 750 3722 755
rect 51 745 60 750
rect 51 740 3722 745
rect 51 735 60 740
rect 51 730 3722 735
rect 51 725 60 730
rect 51 720 3722 725
rect 51 715 60 720
rect 51 710 3722 715
rect 51 705 60 710
rect 51 700 3722 705
rect 51 695 60 700
rect 51 690 3722 695
rect 51 685 60 690
rect 51 680 3722 685
rect 51 675 60 680
rect 51 670 3722 675
rect 51 665 60 670
rect 51 660 3722 665
rect 51 655 60 660
rect 51 650 3722 655
rect 51 645 60 650
rect 51 640 3722 645
rect 51 635 60 640
rect 51 630 3722 635
rect 51 625 60 630
rect 51 620 3722 625
rect 51 615 60 620
rect 51 610 3722 615
rect 51 605 60 610
rect 51 600 3722 605
rect 51 595 60 600
rect 51 590 3722 595
rect 51 585 60 590
rect 51 580 3722 585
rect 51 575 60 580
rect 51 570 3722 575
rect 51 565 60 570
rect 51 560 3722 565
rect 51 555 60 560
rect 51 550 3722 555
rect 51 545 60 550
rect 51 540 3722 545
rect 51 535 60 540
rect 51 530 3722 535
rect 51 525 60 530
rect 51 520 3722 525
rect 51 515 60 520
rect 51 510 3722 515
rect 51 505 60 510
rect 51 500 3722 505
rect 51 495 60 500
rect 51 490 3722 495
rect 51 485 60 490
rect 51 480 3722 485
rect 51 475 60 480
rect 51 470 3722 475
rect 51 465 60 470
rect 51 460 3722 465
rect 51 455 60 460
rect 51 450 3722 455
rect 51 445 60 450
rect 51 440 3722 445
rect 51 435 60 440
rect 51 430 3722 435
rect 51 425 60 430
rect 51 420 3722 425
rect 51 415 60 420
rect 51 410 3722 415
rect 51 405 60 410
rect 51 400 3722 405
rect 51 395 60 400
rect 51 390 3722 395
rect 51 385 60 390
rect 51 380 3722 385
rect 51 375 60 380
rect 51 370 3722 375
rect 51 365 60 370
rect 51 360 3722 365
rect 51 355 60 360
rect 51 350 3722 355
rect 51 345 60 350
rect 51 340 3722 345
rect 51 335 60 340
rect 51 330 3722 335
rect 51 325 60 330
rect 51 320 3722 325
rect 51 315 60 320
rect 51 310 3722 315
rect 51 305 60 310
rect 51 300 3722 305
rect 51 295 60 300
rect 51 290 3722 295
rect 51 285 60 290
rect 51 280 3722 285
rect 51 275 60 280
rect 51 270 3722 275
rect 51 265 60 270
rect 51 260 3722 265
rect 51 255 60 260
rect 51 250 3722 255
rect 51 245 60 250
rect 51 240 3722 245
rect 51 235 60 240
rect 51 230 3722 235
rect 51 225 60 230
rect 51 220 3722 225
rect 51 215 60 220
rect 51 210 3722 215
rect 51 205 60 210
rect 51 200 3722 205
rect 51 195 60 200
rect 51 190 3722 195
rect 51 185 60 190
rect 51 180 3722 185
rect 51 175 60 180
rect 51 170 3722 175
rect 51 165 60 170
rect 51 160 3722 165
rect 51 155 60 160
rect 51 150 3722 155
rect 51 145 60 150
rect 51 140 3722 145
rect 51 135 60 140
rect 51 130 3722 135
rect 51 125 60 130
rect 51 120 3722 125
rect 51 115 60 120
rect 51 110 3722 115
rect 51 105 60 110
rect 51 100 3722 105
rect 51 95 60 100
rect 51 90 3722 95
rect 51 85 60 90
rect 51 80 3722 85
rect 51 75 60 80
rect 51 70 3722 75
rect 51 65 60 70
rect 51 60 3722 65
<< metal3 >>
rect 40 60 46 857
rect 51 855 60 857
rect 51 850 3722 855
rect 51 845 60 850
rect 51 840 3722 845
rect 51 835 60 840
rect 51 830 3722 835
rect 51 825 60 830
rect 51 820 3722 825
rect 51 815 60 820
rect 51 810 3722 815
rect 51 805 60 810
rect 51 800 3722 805
rect 51 795 60 800
rect 51 790 3722 795
rect 51 785 60 790
rect 51 780 3722 785
rect 51 775 60 780
rect 51 770 3722 775
rect 51 765 60 770
rect 51 760 3722 765
rect 51 755 60 760
rect 51 750 3722 755
rect 51 745 60 750
rect 51 740 3722 745
rect 51 735 60 740
rect 51 730 3722 735
rect 51 725 60 730
rect 51 720 3722 725
rect 51 715 60 720
rect 51 710 3722 715
rect 51 705 60 710
rect 51 700 3722 705
rect 51 695 60 700
rect 51 690 3722 695
rect 51 685 60 690
rect 51 680 3722 685
rect 51 675 60 680
rect 51 670 3722 675
rect 51 665 60 670
rect 51 660 3722 665
rect 51 655 60 660
rect 51 650 3722 655
rect 51 645 60 650
rect 51 640 3722 645
rect 51 635 60 640
rect 51 630 3722 635
rect 51 625 60 630
rect 51 620 3722 625
rect 51 615 60 620
rect 51 610 3722 615
rect 51 605 60 610
rect 51 600 3722 605
rect 51 595 60 600
rect 51 590 3722 595
rect 51 585 60 590
rect 51 580 3722 585
rect 51 575 60 580
rect 51 570 3722 575
rect 51 565 60 570
rect 51 560 3722 565
rect 51 555 60 560
rect 51 550 3722 555
rect 51 545 60 550
rect 51 540 3722 545
rect 51 535 60 540
rect 51 530 3722 535
rect 51 525 60 530
rect 51 520 3722 525
rect 51 515 60 520
rect 51 510 3722 515
rect 51 505 60 510
rect 51 500 3722 505
rect 51 495 60 500
rect 51 490 3722 495
rect 51 485 60 490
rect 51 480 3722 485
rect 51 475 60 480
rect 51 470 3722 475
rect 51 465 60 470
rect 51 460 3722 465
rect 51 455 60 460
rect 51 450 3722 455
rect 51 445 60 450
rect 51 440 3722 445
rect 51 435 60 440
rect 51 430 3722 435
rect 51 425 60 430
rect 51 420 3722 425
rect 51 415 60 420
rect 51 410 3722 415
rect 51 405 60 410
rect 51 400 3722 405
rect 51 395 60 400
rect 51 390 3722 395
rect 51 385 60 390
rect 51 380 3722 385
rect 51 375 60 380
rect 51 370 3722 375
rect 51 365 60 370
rect 51 360 3722 365
rect 51 355 60 360
rect 51 350 3722 355
rect 51 345 60 350
rect 51 340 3722 345
rect 51 335 60 340
rect 51 330 3722 335
rect 51 325 60 330
rect 51 320 3722 325
rect 51 315 60 320
rect 51 310 3722 315
rect 51 305 60 310
rect 51 300 3722 305
rect 51 295 60 300
rect 51 290 3722 295
rect 51 285 60 290
rect 51 280 3722 285
rect 51 275 60 280
rect 51 270 3722 275
rect 51 265 60 270
rect 51 260 3722 265
rect 51 255 60 260
rect 51 250 3722 255
rect 51 245 60 250
rect 51 240 3722 245
rect 51 235 60 240
rect 51 230 3722 235
rect 51 225 60 230
rect 51 220 3722 225
rect 51 215 60 220
rect 51 210 3722 215
rect 51 205 60 210
rect 51 200 3722 205
rect 51 195 60 200
rect 51 190 3722 195
rect 51 185 60 190
rect 51 180 3722 185
rect 51 175 60 180
rect 51 170 3722 175
rect 51 165 60 170
rect 51 160 3722 165
rect 51 155 60 160
rect 51 150 3722 155
rect 51 145 60 150
rect 51 140 3722 145
rect 51 135 60 140
rect 51 130 3722 135
rect 51 125 60 130
rect 51 120 3722 125
rect 51 115 60 120
rect 51 110 3722 115
rect 51 105 60 110
rect 51 100 3722 105
rect 51 95 60 100
rect 51 90 3722 95
rect 51 85 60 90
rect 51 80 3722 85
rect 51 75 60 80
rect 51 70 3722 75
rect 51 65 60 70
rect 51 60 3722 65
<< m234contact >>
rect 20 429 28 497
rect 46 60 51 857
<< metal4 >>
rect 19 429 20 497
rect 40 60 46 857
rect 51 60 52 857
rect 60 850 3722 855
rect 60 840 3722 845
rect 60 830 3722 835
rect 60 820 3722 825
rect 60 810 3722 815
rect 60 800 3722 805
rect 60 790 3722 795
rect 60 780 3722 785
rect 60 770 3722 775
rect 60 760 3722 765
rect 60 750 3722 755
rect 60 740 3722 745
rect 60 730 3722 735
rect 60 720 3722 725
rect 60 710 3722 715
rect 60 700 3722 705
rect 60 690 3722 695
rect 60 680 3722 685
rect 60 670 3722 675
rect 60 660 3722 665
rect 60 650 3722 655
rect 60 640 3722 645
rect 60 630 3722 635
rect 60 620 3722 625
rect 60 610 3722 615
rect 60 600 3722 605
rect 60 590 3722 595
rect 60 580 3722 585
rect 60 570 3722 575
rect 60 560 3722 565
rect 60 550 3722 555
rect 60 540 3722 545
rect 60 530 3722 535
rect 60 520 3722 525
rect 60 510 3722 515
rect 60 500 3722 505
rect 60 490 3722 495
rect 60 480 3722 485
rect 60 470 3722 475
rect 60 460 3722 465
rect 60 450 3722 455
rect 60 440 3722 445
rect 60 430 3722 435
rect 60 420 3722 425
rect 60 410 3722 415
rect 60 400 3722 405
rect 60 390 3722 395
rect 60 380 3722 385
rect 60 370 3722 375
rect 60 360 3722 365
rect 60 350 3722 355
rect 60 340 3722 345
rect 60 330 3722 335
rect 60 320 3722 325
rect 60 310 3722 315
rect 60 300 3722 305
rect 60 290 3722 295
rect 60 280 3722 285
rect 60 270 3722 275
rect 60 260 3722 265
rect 60 250 3722 255
rect 60 240 3722 245
rect 60 230 3722 235
rect 60 220 3722 225
rect 60 210 3722 215
rect 60 200 3722 205
rect 60 190 3722 195
rect 60 180 3722 185
rect 60 170 3722 175
rect 60 160 3722 165
rect 60 150 3722 155
rect 60 140 3722 145
rect 60 130 3722 135
rect 60 120 3722 125
rect 60 110 3722 115
rect 60 100 3722 105
rect 60 90 3722 95
rect 60 80 3722 85
rect 60 70 3722 75
rect 60 60 3722 65
<< metal5 >>
rect 40 60 52 857
rect 60 850 3722 855
rect 60 840 3722 845
rect 60 830 3722 835
rect 60 820 3722 825
rect 60 810 3722 815
rect 60 800 3722 805
rect 60 790 3722 795
rect 60 780 3722 785
rect 60 770 3722 775
rect 60 760 3722 765
rect 60 750 3722 755
rect 60 740 3722 745
rect 60 730 3722 735
rect 60 720 3722 725
rect 60 710 3722 715
rect 60 700 3722 705
rect 60 690 3722 695
rect 60 680 3722 685
rect 60 670 3722 675
rect 60 660 3722 665
rect 60 650 3722 655
rect 60 640 3722 645
rect 60 630 3722 635
rect 60 620 3722 625
rect 60 610 3722 615
rect 60 600 3722 605
rect 60 590 3722 595
rect 60 580 3722 585
rect 60 570 3722 575
rect 60 560 3722 565
rect 60 550 3722 555
rect 60 540 3722 545
rect 60 530 3722 535
rect 60 520 3722 525
rect 60 510 3722 515
rect 60 500 3722 505
rect 60 490 3722 495
rect 60 480 3722 485
rect 60 470 3722 475
rect 60 460 3722 465
rect 60 450 3722 455
rect 60 440 3722 445
rect 60 430 3722 435
rect 60 420 3722 425
rect 60 410 3722 415
rect 60 400 3722 405
rect 60 390 3722 395
rect 60 380 3722 385
rect 60 370 3722 375
rect 60 360 3722 365
rect 60 350 3722 355
rect 60 340 3722 345
rect 60 330 3722 335
rect 60 320 3722 325
rect 60 310 3722 315
rect 60 300 3722 305
rect 60 290 3722 295
rect 60 280 3722 285
rect 60 270 3722 275
rect 60 260 3722 265
rect 60 250 3722 255
rect 60 240 3722 245
rect 60 230 3722 235
rect 60 220 3722 225
rect 60 210 3722 215
rect 60 200 3722 205
rect 60 190 3722 195
rect 60 180 3722 185
rect 60 170 3722 175
rect 60 160 3722 165
rect 60 150 3722 155
rect 60 140 3722 145
rect 60 130 3722 135
rect 60 120 3722 125
rect 60 110 3722 115
rect 60 100 3722 105
rect 60 90 3722 95
rect 60 80 3722 85
rect 60 70 3722 75
rect 60 60 3722 65
<< m456contact >>
rect 11 429 19 497
rect 52 60 60 857
<< metal6 >>
rect -52 429 11 497
rect 40 60 52 857
rect 60 850 3722 855
rect 60 840 3722 845
rect 60 830 3722 835
rect 60 820 3722 825
rect 60 810 3722 815
rect 60 800 3722 805
rect 60 790 3722 795
rect 60 780 3722 785
rect 60 770 3722 775
rect 60 760 3722 765
rect 60 750 3722 755
rect 60 740 3722 745
rect 60 730 3722 735
rect 60 720 3722 725
rect 60 710 3722 715
rect 60 700 3722 705
rect 60 690 3722 695
rect 60 680 3722 685
rect 60 670 3722 675
rect 60 660 3722 665
rect 60 650 3722 655
rect 60 640 3722 645
rect 60 630 3722 635
rect 60 620 3722 625
rect 60 610 3722 615
rect 60 600 3722 605
rect 60 590 3722 595
rect 60 580 3722 585
rect 60 570 3722 575
rect 60 560 3722 565
rect 60 550 3722 555
rect 60 540 3722 545
rect 60 530 3722 535
rect 60 520 3722 525
rect 60 510 3722 515
rect 60 500 3722 505
rect 60 490 3722 495
rect 60 480 3722 485
rect 60 470 3722 475
rect 60 460 3722 465
rect 60 450 3722 455
rect 60 440 3722 445
rect 60 430 3722 435
rect 60 420 3722 425
rect 60 410 3722 415
rect 60 400 3722 405
rect 60 390 3722 395
rect 60 380 3722 385
rect 60 370 3722 375
rect 60 360 3722 365
rect 60 350 3722 355
rect 60 340 3722 345
rect 60 330 3722 335
rect 60 320 3722 325
rect 60 310 3722 315
rect 60 300 3722 305
rect 60 290 3722 295
rect 60 280 3722 285
rect 60 270 3722 275
rect 60 260 3722 265
rect 60 250 3722 255
rect 60 240 3722 245
rect 60 230 3722 235
rect 60 220 3722 225
rect 60 210 3722 215
rect 60 200 3722 205
rect 60 190 3722 195
rect 60 180 3722 185
rect 60 170 3722 175
rect 60 160 3722 165
rect 60 150 3722 155
rect 60 140 3722 145
rect 60 130 3722 135
rect 60 120 3722 125
rect 60 110 3722 115
rect 60 100 3722 105
rect 60 90 3722 95
rect 60 80 3722 85
rect 60 70 3722 75
rect 60 60 3722 65
<< labels >>
rlabel metal6 -20 463 -20 463 1 ninepF
<< end >>
