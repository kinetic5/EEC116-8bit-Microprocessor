magic
tech scmos
timestamp 1575407437
<< ntransistor >>
rect 10 28 12 32
rect 30 28 32 32
rect 40 28 42 32
rect 60 28 62 32
<< ptransistor >>
rect 10 44 12 50
rect 30 44 32 50
rect 40 44 42 50
rect 60 44 62 50
<< ndiffusion >>
rect 9 28 10 32
rect 12 28 13 32
rect 29 28 30 32
rect 32 28 33 32
rect 39 28 40 32
rect 42 28 43 32
rect 59 28 60 32
rect 62 28 63 32
<< pdiffusion >>
rect 6 48 10 50
rect 9 44 10 48
rect 12 48 16 50
rect 12 44 13 48
rect 26 48 30 50
rect 29 44 30 48
rect 32 48 40 50
rect 32 44 33 48
rect 39 44 40 48
rect 42 48 46 50
rect 42 44 43 48
rect 56 49 60 50
rect 59 44 60 49
rect 62 48 66 50
rect 62 44 63 48
<< ndcontact >>
rect 3 28 9 32
rect 13 28 19 32
rect 23 28 29 32
rect 33 28 39 32
rect 43 28 48 32
rect 53 28 59 32
rect 63 28 69 32
<< pdcontact >>
rect 3 44 9 48
rect 13 44 19 48
rect 23 44 29 48
rect 33 44 39 48
rect 43 44 48 48
rect 63 44 69 48
<< polysilicon >>
rect 0 20 2 56
rect 10 50 12 56
rect 10 41 12 44
rect 10 32 12 36
rect 10 20 12 28
rect 20 20 22 56
rect 30 50 32 51
rect 40 50 42 52
rect 30 41 32 44
rect 40 41 42 44
rect 30 32 32 35
rect 40 32 42 35
rect 30 25 32 28
rect 40 25 42 28
rect 40 20 42 21
rect 50 20 52 55
rect 60 50 62 52
rect 60 40 62 44
rect 60 32 62 35
rect 60 20 62 28
rect 70 20 72 56
rect 80 20 82 56
rect 90 20 92 56
rect 100 20 102 56
rect 110 20 112 56
rect 120 20 122 56
rect 130 20 132 56
rect 140 20 142 56
rect 150 20 152 56
rect 160 20 162 56
<< polycontact >>
rect 40 52 44 56
rect 40 21 44 25
rect 58 52 62 56
<< metal1 >>
rect 0 66 122 74
rect 3 48 9 66
rect 40 56 62 57
rect 44 53 58 56
rect 19 44 23 48
rect 23 32 29 44
rect 19 28 23 32
rect 33 38 39 44
rect 33 33 34 38
rect 33 32 39 33
rect 43 41 48 44
rect 43 32 48 36
rect 52 44 54 49
rect 65 48 70 66
rect 69 44 70 48
rect 52 32 56 44
rect 52 28 53 32
rect 69 28 70 32
rect 3 10 9 28
rect 52 25 56 28
rect 44 21 56 25
rect 65 10 70 28
rect 0 2 122 10
<< m2contact >>
rect 34 33 39 38
rect 43 36 48 41
<< pm12contact >>
rect 30 51 35 56
rect 9 36 14 41
rect 59 35 64 40
rect 29 20 34 25
<< pdm12contact >>
rect 54 44 59 49
<< metal2 >>
rect 54 49 59 51
rect 9 41 14 42
rect 43 41 48 42
rect 59 25 64 35
<< m3contact >>
rect 35 51 40 56
rect 54 51 59 56
rect 9 42 14 47
rect 43 42 48 47
rect 34 20 39 25
rect 59 20 64 25
<< metal3 >>
rect 40 51 54 56
rect 14 42 43 47
rect 39 20 59 25
<< labels >>
rlabel metal1 3 70 3 70 4 Vdd
rlabel metal1 3 6 3 6 2 Gnd
rlabel m2contact 36 35 36 35 1 z
rlabel pm12contact 61 38 61 38 1 a
rlabel pm12contact 11 38 11 38 1 b
<< end >>
