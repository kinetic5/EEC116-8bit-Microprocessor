magic
tech scmos
timestamp 1575763138
<< ntransistor >>
rect -96 -13 -94 -9
rect -86 -13 -84 -9
rect -66 -13 -64 -9
rect -56 -13 -54 -9
rect -46 -21 -44 -17
rect -26 -13 -24 -9
rect -16 -13 -14 -9
rect -6 -13 -4 -9
rect 4 -13 6 -9
rect 14 -21 16 -17
rect 34 -13 36 -9
rect 44 -13 46 -9
rect 54 -21 56 -17
<< ptransistor >>
rect -46 20 -44 25
rect -96 11 -94 17
rect -86 11 -84 17
rect -66 11 -64 17
rect -56 11 -54 17
rect 14 20 16 25
rect -26 11 -24 17
rect -16 11 -14 17
rect -6 11 -4 17
rect 4 11 6 17
rect 54 20 56 25
rect 34 11 36 17
rect 44 11 46 17
<< ndiffusion >>
rect -97 -13 -96 -9
rect -94 -13 -93 -9
rect -87 -13 -86 -9
rect -84 -13 -83 -9
rect -67 -13 -66 -9
rect -64 -13 -62 -9
rect -58 -13 -56 -9
rect -54 -13 -53 -9
rect -52 -21 -46 -17
rect -44 -21 -41 -17
rect -32 -13 -31 -9
rect -27 -13 -26 -9
rect -24 -13 -22 -9
rect -17 -13 -16 -9
rect -14 -13 -12 -9
rect -8 -13 -6 -9
rect -4 -13 -3 -9
rect 3 -13 4 -9
rect 6 -13 8 -9
rect 9 -21 14 -17
rect 16 -21 18 -17
rect 32 -13 34 -9
rect 36 -13 37 -9
rect 43 -13 44 -9
rect 46 -13 48 -9
rect 53 -21 54 -17
rect 56 -21 58 -17
rect -51 -24 -47 -21
rect 9 -24 13 -21
<< pdiffusion >>
rect -51 25 -47 29
rect 9 25 13 28
rect -51 20 -46 25
rect -44 20 -42 25
rect -97 11 -96 17
rect -94 11 -93 17
rect -87 11 -86 17
rect -84 11 -83 17
rect -72 16 -66 17
rect -67 11 -66 16
rect -64 11 -62 17
rect -58 11 -56 17
rect -54 16 -48 17
rect -54 11 -52 16
rect 9 20 14 25
rect 16 20 18 25
rect -32 11 -31 17
rect -27 11 -26 17
rect -24 11 -23 17
rect -17 11 -16 17
rect -14 11 -13 17
rect -7 11 -6 17
rect -4 11 -3 17
rect 3 11 4 17
rect 6 16 12 17
rect 6 11 8 16
rect 53 21 54 25
rect 48 20 54 21
rect 56 20 58 25
rect 32 11 34 17
rect 36 11 37 17
rect 43 11 44 17
rect 46 16 52 17
rect 46 11 48 16
<< ndcontact >>
rect -102 -13 -97 -9
rect -93 -13 -87 -9
rect -83 -13 -78 -9
rect -73 -13 -67 -9
rect -62 -13 -58 -9
rect -53 -13 -49 -9
rect -41 -21 -37 -17
rect -31 -13 -27 -9
rect -22 -13 -17 -9
rect -12 -13 -8 -9
rect -3 -13 3 -9
rect 8 -13 12 -9
rect 18 -21 22 -17
rect 28 -13 32 -9
rect 37 -13 43 -9
rect 48 -13 52 -9
rect 48 -21 53 -17
rect 58 -21 62 -17
rect -51 -28 -47 -24
rect 9 -28 13 -24
<< pdcontact >>
rect -51 29 -47 33
rect 9 28 13 32
rect -42 20 -38 25
rect -102 11 -97 17
rect -93 11 -87 17
rect -83 11 -78 17
rect -62 11 -58 17
rect -52 11 -48 16
rect 18 20 22 25
rect -31 11 -27 17
rect -23 11 -17 17
rect -13 11 -7 17
rect -3 11 3 17
rect 8 11 12 16
rect 48 21 53 25
rect 58 20 62 25
rect 28 11 32 17
rect 37 11 43 17
rect 48 11 52 16
<< psubstratepcontact >>
rect -65 -30 -57 -24
rect -23 -31 -11 -24
rect 27 -31 43 -24
<< nsubstratencontact >>
rect -64 29 -55 35
rect -26 28 -11 35
rect 26 28 42 35
<< polysilicon >>
rect -46 25 -44 28
rect 14 25 16 28
rect 54 25 56 28
rect -106 -16 -104 20
rect -96 17 -94 20
rect -86 17 -84 20
rect -96 -1 -94 11
rect -86 8 -84 11
rect -96 -9 -94 -6
rect -86 -9 -84 3
rect -96 -16 -94 -13
rect -86 -16 -84 -13
rect -76 -16 -74 20
rect -66 17 -64 20
rect -56 17 -54 20
rect -66 4 -64 11
rect -56 4 -54 11
rect -46 -1 -44 20
rect -66 -9 -64 -2
rect -56 -9 -54 -2
rect -66 -16 -64 -13
rect -56 -16 -54 -13
rect -46 -17 -44 -6
rect -36 -21 -34 25
rect -26 17 -24 25
rect -16 17 -14 25
rect -6 17 -4 20
rect 4 17 6 20
rect -26 -9 -24 11
rect -16 -1 -14 11
rect -6 4 -4 11
rect 4 4 6 11
rect 14 -1 16 20
rect -16 -9 -14 -6
rect -6 -9 -4 -2
rect 4 -9 6 -2
rect -26 -16 -24 -13
rect -16 -21 -14 -13
rect -6 -16 -4 -13
rect 4 -16 6 -13
rect 14 -17 16 -6
rect 24 -21 26 25
rect 34 17 36 25
rect 44 17 46 25
rect 34 -1 36 11
rect 44 -1 46 11
rect 54 -1 56 20
rect 34 -9 36 -6
rect 44 -9 46 -6
rect 34 -21 36 -13
rect 44 -21 46 -13
rect 54 -17 56 -6
rect 64 -21 66 25
rect -46 -24 -44 -21
rect 14 -24 16 -21
rect 54 -24 56 -21
<< polycontact >>
rect -96 -6 -92 -1
rect 43 -6 47 -1
<< metal1 >>
rect -108 35 68 36
rect -108 29 -64 35
rect -55 33 -26 35
rect -55 29 -51 33
rect -47 29 -26 33
rect -108 28 -26 29
rect -11 32 26 35
rect -11 28 9 32
rect 13 28 26 32
rect 42 28 68 35
rect -91 17 -87 28
rect -103 11 -102 17
rect -78 11 -76 17
rect -103 -9 -99 6
rect -80 -9 -76 11
rect -103 -13 -102 -9
rect -78 -13 -76 -9
rect -73 11 -72 16
rect -73 -9 -68 11
rect -62 -2 -58 11
rect -53 11 -52 16
rect -53 8 -50 11
rect -62 -7 -61 -2
rect -62 -9 -58 -7
rect -53 -9 -50 3
rect -93 -24 -87 -13
rect -38 -17 -34 25
rect -23 17 -17 28
rect 22 20 23 25
rect -31 8 -27 11
rect -31 -9 -27 3
rect -10 -9 -7 11
rect -17 -13 -16 -9
rect -8 -13 -7 -9
rect -3 0 3 11
rect -3 -6 -2 0
rect -3 -9 3 -6
rect 6 11 8 16
rect 6 10 12 11
rect 6 5 8 10
rect 6 -9 9 5
rect 6 -13 8 -9
rect 20 -10 23 20
rect 37 17 43 28
rect 48 25 53 28
rect 62 20 63 25
rect 52 11 54 16
rect 28 10 31 11
rect 28 -9 31 5
rect 50 -1 54 11
rect 39 -6 43 -1
rect 50 -6 51 -1
rect 50 -9 54 -6
rect -37 -21 -28 -17
rect -20 -24 -16 -13
rect 52 -13 54 -9
rect 19 -17 23 -15
rect 22 -21 23 -17
rect 37 -24 43 -13
rect 59 -17 63 20
rect 62 -21 63 -17
rect 48 -24 53 -21
rect -108 -30 -65 -24
rect -57 -28 -51 -24
rect -47 -28 -23 -24
rect -57 -30 -23 -28
rect -108 -31 -23 -30
rect -11 -28 9 -24
rect 13 -28 27 -24
rect -11 -31 27 -28
rect 43 -31 68 -24
rect -108 -32 68 -31
<< m2contact >>
rect -92 -6 -87 -1
rect -53 3 -48 8
rect -61 -7 -56 -2
rect -81 -18 -76 -13
rect -31 3 -26 8
rect -2 -6 3 0
rect 8 5 13 10
rect 26 5 31 10
rect 19 -15 24 -10
<< pm12contact >>
rect -68 20 -63 25
rect -58 20 -53 25
rect -88 3 -83 8
rect -47 -6 -42 -1
rect -68 -21 -63 -16
rect -58 -21 -53 -16
rect -8 20 -3 25
rect 2 20 7 25
rect -18 -6 -13 -1
rect 12 -6 17 -1
rect 34 -6 39 -1
rect 51 -6 56 -1
rect -28 -21 -23 -16
rect -8 -21 -3 -16
rect 2 -21 7 -16
<< pdm12contact >>
rect -72 11 -67 16
<< metal2 >>
rect -69 30 6 33
rect -64 29 6 30
rect 1 25 6 29
rect -59 20 -58 25
rect -53 20 -13 25
rect 1 20 2 25
rect -59 16 -56 20
rect -62 13 -56 16
rect 1 17 6 20
rect -62 6 -58 13
rect 1 9 4 17
rect -70 2 -58 6
rect -48 3 -31 8
rect -9 5 4 9
rect 13 5 26 10
rect -92 -13 -87 -6
rect -70 -13 -66 2
rect -56 -6 -47 -2
rect -56 -7 -42 -6
rect -28 -6 -18 -3
rect -28 -7 -14 -6
rect -92 -18 -81 -13
rect -76 -16 -66 -13
rect -28 -16 -23 -7
rect -76 -18 -68 -16
rect -70 -21 -68 -18
rect -9 -16 -6 5
rect 3 -6 12 -1
rect 34 -10 38 -6
rect 24 -15 38 -10
rect -9 -21 -8 -16
<< m3contact >>
rect -69 25 -64 30
rect -13 20 -8 25
rect -53 -21 -48 -16
rect 7 -21 12 -16
<< m123contact >>
rect -103 6 -97 11
<< metal3 >>
rect -103 25 -69 29
rect -103 23 -64 25
rect -103 11 -97 23
rect -69 -16 -64 23
rect -8 20 -3 25
rect -8 9 -4 20
rect -8 4 6 9
rect 1 -16 6 4
rect -69 -21 -53 -16
rect 1 -21 7 -16
<< labels >>
rlabel metal1 12 32 12 32 1 Vdd
rlabel metal1 0 -30 0 -30 1 Gnd
rlabel metal1 -71 1 -71 1 1 D
rlabel pm12contact -86 5 -86 5 1 clk
rlabel metal1 61 6 61 6 1 Qbar
rlabel pm12contact 54 -4 54 -4 1 Q
<< end >>
