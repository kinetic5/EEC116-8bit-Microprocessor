magic
tech scmos
timestamp 1575836395
<< error_s >>
rect -194 85 -193 86
rect 46 85 47 86
rect 286 85 287 86
rect 526 85 527 86
rect 766 85 767 86
rect 1006 85 1007 86
rect 1246 85 1247 86
rect 1486 85 1487 86
<< metal1 >>
rect 1674 133 1785 141
rect 1679 74 1687 82
rect 1695 74 1764 82
rect 1777 70 1785 133
rect 1679 62 1687 70
rect 1695 62 1785 70
<< metal2 >>
rect -43 154 1657 159
rect -28 109 -23 154
rect 212 114 217 154
rect 452 109 457 154
rect 692 109 697 154
rect 932 109 937 154
rect 1172 109 1177 154
rect 1412 109 1417 154
rect 1652 109 1657 154
rect -184 67 -178 72
rect 56 -6 62 0
rect 296 -78 302 -72
rect 536 -150 542 -144
rect 776 -222 782 -216
rect 1016 -295 1022 -288
rect 1256 -366 1262 -360
rect 1496 -437 1502 -432
<< m123contact >>
rect 1687 74 1695 82
rect 1687 62 1695 70
<< metal3 >>
rect -38 141 -32 151
rect 202 137 208 149
rect 442 137 448 149
rect 682 137 688 150
rect 922 137 928 150
rect 1162 137 1168 150
rect 1402 137 1408 150
rect 1642 137 1648 153
rect 231 -8 239 0
rect 471 -80 479 -72
rect 711 -152 719 -144
rect 951 -224 959 -216
rect 1191 -296 1199 -288
rect 1431 -368 1439 -360
<< m345contact >>
rect 1695 74 1703 82
rect 1695 62 1703 70
<< metal5 >>
rect -249 123 -241 130
rect -9 51 -1 58
rect 231 -21 239 -14
rect 471 -93 479 -86
rect 711 -165 719 -158
rect 951 -237 959 -230
rect 1191 -309 1199 -302
rect 1431 -381 1439 -374
<< m6contact >>
rect 1703 75 1711 83
rect 1703 62 1711 70
<< metal6 >>
rect 1633 -370 1641 156
rect 1649 84 1657 156
rect 1649 83 1711 84
rect 1649 76 1703 83
rect 1649 -430 1657 76
use mult_and  mult_and_0
array 0 7 240 0 0 72
timestamp 1575836395
transform 1 0 -488 0 1 64
box 247 8 487 78
use mult_hadder  mult_hadder_0
timestamp 1575779281
transform 1 0 -7 0 1 -7
box 6 7 246 79
use mult_fadder  mult_fadder_0
array 0 5 240 0 0 72
timestamp 1575623072
transform 1 0 233 0 1 -8
box 6 8 246 80
use mult_hadder  mult_hadder_1
timestamp 1575779281
transform 1 0 233 0 1 -79
box 6 7 246 79
use mult_fadder  mult_fadder_1
array 0 4 240 0 0 72
timestamp 1575623072
transform 1 0 473 0 1 -80
box 6 8 246 80
use mult_hadder  mult_hadder_2
timestamp 1575779281
transform 1 0 473 0 1 -151
box 6 7 246 79
use mult_fadder  mult_fadder_2
array 0 3 240 0 0 72
timestamp 1575623072
transform 1 0 713 0 1 -152
box 6 8 246 80
use mult_hadder  mult_hadder_3
timestamp 1575779281
transform 1 0 713 0 1 -223
box 6 7 246 79
use mult_fadder  mult_fadder_3
array 0 2 240 0 0 72
timestamp 1575623072
transform 1 0 953 0 1 -224
box 6 8 246 80
use mult_hadder  mult_hadder_4
timestamp 1575779281
transform 1 0 953 0 1 -295
box 6 7 246 79
use mult_fadder  mult_fadder_4
array 0 1 240 0 0 72
timestamp 1575623072
transform 1 0 1193 0 1 -296
box 6 8 246 80
use mult_hadder  mult_hadder_5
timestamp 1575779281
transform 1 0 1193 0 1 -367
box 6 7 246 79
use mult_fadder  mult_fadder_5
timestamp 1575623072
transform 1 0 1433 0 1 -368
box 6 8 246 80
use mult_hadder  mult_hadder_6
timestamp 1575779281
transform 1 0 1433 0 1 -439
box 6 7 246 79
<< labels >>
rlabel metal5 -5 54 -5 54 3 y1
rlabel metal5 235 -17 235 -17 1 y2
rlabel metal5 475 -90 475 -90 1 y3
rlabel metal5 715 -161 715 -161 1 y4
rlabel metal5 955 -233 955 -233 1 y5
rlabel metal5 1195 -306 1195 -306 1 y6
rlabel metal5 1435 -377 1435 -377 1 y7
rlabel metal2 59 -3 59 -3 1 z1
rlabel metal2 299 -75 299 -75 1 z2
rlabel metal2 539 -147 539 -147 1 z3
rlabel metal2 779 -219 779 -219 1 z4
rlabel metal2 1019 -291 1019 -291 1 z5
rlabel metal2 1259 -364 1259 -364 1 z6
rlabel metal2 1499 -434 1499 -434 1 z7
rlabel metal2 -181 71 -181 71 1 z0
rlabel metal5 -245 126 -245 126 3 y0
rlabel metal6 1653 78 1653 78 5 Gnd
rlabel metal6 1637 78 1637 78 5 Vdd
rlabel metal2 -25 156 -25 156 5 clk
rlabel metal3 -35 147 -35 147 1 x0
rlabel metal3 205 146 205 146 1 x1
rlabel metal3 444 146 444 146 1 x2
rlabel metal3 685 146 685 146 1 x3
rlabel metal3 925 147 925 147 1 x4
rlabel metal3 1165 147 1165 147 1 x5
rlabel metal3 1645 147 1645 147 1 x7
rlabel metal3 1405 147 1405 147 1 x6
<< end >>
