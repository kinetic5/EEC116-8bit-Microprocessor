magic
tech scmos
timestamp 1575772227
<< ntransistor >>
rect 10 25 12 29
rect 20 25 22 29
rect 30 23 32 29
<< ptransistor >>
rect 10 45 12 51
rect 30 50 32 59
rect 20 41 22 47
<< ndiffusion >>
rect 9 25 10 29
rect 12 25 13 29
rect 19 25 20 29
rect 22 25 23 29
rect 29 23 30 29
rect 32 23 33 29
<< pdiffusion >>
rect 9 45 10 51
rect 12 47 18 51
rect 29 51 30 59
rect 26 50 30 51
rect 32 56 39 59
rect 32 50 33 56
rect 12 45 20 47
rect 13 41 20 45
rect 22 46 26 47
rect 22 41 23 46
<< ndcontact >>
rect 3 25 9 29
rect 13 25 19 29
rect 23 23 29 29
rect 33 23 39 29
<< pdcontact >>
rect 3 45 9 51
rect 23 51 29 59
rect 23 41 29 46
<< polysilicon >>
rect 0 14 2 62
rect 10 51 12 62
rect 20 47 22 62
rect 30 59 32 62
rect 10 38 12 45
rect 20 38 22 41
rect 30 39 32 50
rect 10 29 12 32
rect 20 29 22 32
rect 30 29 32 33
rect 10 14 12 25
rect 20 14 22 25
rect 30 14 32 23
rect 40 14 42 62
<< metal1 >>
rect 0 64 42 72
rect 3 51 9 64
rect 23 59 29 64
rect 39 50 40 56
rect 29 41 32 46
rect 26 39 32 41
rect 26 33 28 39
rect 36 29 40 50
rect 3 12 9 25
rect 39 23 40 29
rect 23 12 29 23
rect 0 4 42 12
<< m2contact >>
rect 13 19 19 25
<< pm12contact >>
rect 8 32 13 38
rect 18 32 23 38
rect 28 33 33 39
<< pdm12contact >>
rect 33 50 39 56
<< metal2 >>
rect 27 33 28 39
rect 27 28 32 33
rect 13 25 32 28
rect 19 23 32 25
<< m3contact >>
rect 33 44 39 50
rect 7 38 13 44
rect 17 38 23 44
<< metal3 >>
rect 33 23 39 44
<< labels >>
rlabel metal1 3 68 3 68 4 Vdd
rlabel metal1 3 8 3 8 2 Gnd
rlabel m3contact 20 41 20 41 1 or_a
rlabel m3contact 10 41 10 41 1 or_b
rlabel metal3 36 26 36 26 1 or_z
<< end >>
