magic
tech scmos
timestamp 1575532970
<< metal2 >>
rect -136 144 -130 149
rect 96 144 102 149
rect 328 144 334 149
rect 560 144 566 149
rect 792 144 798 149
rect 1024 144 1030 149
rect 1256 144 1262 149
rect 1488 144 1494 149
rect -123 68 -118 72
rect 109 68 114 72
rect 109 -3 114 2
rect 341 -75 346 -70
rect 573 -147 578 -142
rect 805 -219 810 -214
rect 1037 -291 1042 -286
rect 1269 -363 1274 -358
rect 1501 -435 1506 -430
<< metal3 >>
rect -239 127 -232 133
rect -7 65 0 72
rect 1396 70 1401 75
rect -5 56 0 61
rect -6 8 0 46
rect -6 2 12 8
rect 225 -7 232 0
rect 227 -16 232 -11
rect 226 -64 232 -26
rect 226 -70 244 -64
rect 457 -79 464 -72
rect 459 -88 464 -83
rect 458 -136 464 -98
rect 458 -142 476 -136
rect 689 -151 696 -144
rect 691 -160 696 -155
rect 690 -208 696 -170
rect 690 -214 708 -208
rect 921 -223 928 -216
rect 923 -232 928 -227
rect 922 -280 928 -242
rect 922 -286 940 -280
rect 1153 -295 1160 -288
rect 1155 -304 1160 -299
rect 1154 -352 1160 -314
rect 1154 -358 1172 -352
rect 1385 -367 1392 -360
rect 1387 -376 1392 -371
rect 1386 -424 1392 -386
rect 1386 -430 1404 -424
<< metal4 >>
rect 1396 -430 1420 162
rect 1573 -370 1597 164
use pand  pand_0
array 0 7 232 0 0 72
timestamp 1575507270
transform 1 0 -232 0 1 136
box 0 -64 232 8
use psum  psum_0
array 0 6 232 0 0 72
timestamp 1575532930
transform 1 0 40 0 1 -2
box -43 2 195 74
use psum  psum_1
array 0 5 232 0 0 72
timestamp 1575532930
transform 1 0 272 0 1 -74
box -43 2 195 74
use psum  psum_2
array 0 4 232 0 0 72
timestamp 1575532930
transform 1 0 504 0 1 -146
box -43 2 195 74
use psum  psum_3
array 0 3 232 0 0 72
timestamp 1575532930
transform 1 0 736 0 1 -218
box -43 2 195 74
use psum  psum_4
array 0 2 232 0 0 72
timestamp 1575532930
transform 1 0 968 0 1 -290
box -43 2 195 74
use psum  psum_5
array 0 1 232 0 0 72
timestamp 1575532930
transform 1 0 1200 0 1 -362
box -43 2 195 74
use psum  psum_6
timestamp 1575532930
transform 1 0 1432 0 1 -434
box -43 2 195 74
<< labels >>
rlabel metal4 1408 78 1408 78 5 Gnd
rlabel metal4 1585 76 1585 76 1 Vdd
rlabel metal3 -3 58 -3 58 3 y1
rlabel metal3 230 -14 230 -14 1 y2
rlabel metal3 461 -86 461 -86 1 y3
rlabel metal3 693 -157 693 -157 1 y4
rlabel metal3 925 -230 925 -230 1 y5
rlabel metal3 1157 -302 1157 -302 1 y6
rlabel metal3 1389 -374 1389 -374 1 y7
rlabel metal2 112 -1 112 -1 1 z1
rlabel metal2 344 -73 344 -73 1 z2
rlabel metal2 576 -145 576 -145 1 z3
rlabel metal2 807 -217 807 -217 1 z4
rlabel metal2 1039 -288 1039 -288 1 z5
rlabel metal2 1271 -360 1271 -360 1 z6
rlabel metal2 1503 -432 1503 -432 1 z7
rlabel metal3 -236 130 -236 130 3 y0
rlabel metal2 -121 70 -121 70 1 z0
rlabel metal2 -133 146 -133 146 1 x0
rlabel metal2 98 146 98 146 1 x1
rlabel metal2 331 145 331 145 1 x2
rlabel metal2 563 146 563 146 1 x3
rlabel metal2 795 146 795 146 1 x4
rlabel metal2 1027 146 1027 146 1 x5
rlabel metal2 1259 146 1259 146 1 x6
rlabel metal2 1490 146 1490 146 1 x7
rlabel metal2 111 70 111 70 1 z1_p
rlabel metal3 -3 42 -3 42 1 z1_cin
rlabel metal3 -4 68 -4 68 1 z1_x
<< end >>
