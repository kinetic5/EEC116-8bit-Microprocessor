magic
tech scmos
timestamp 1576135017
<< nwell >>
rect -76 -87 134 -50
<< pwell >>
rect -76 -89 134 -87
rect -83 -101 134 -89
rect -76 -122 134 -101
<< ntransistor >>
rect -62 -97 -60 -93
rect -52 -97 -50 -93
rect -42 -97 -40 -93
rect -32 -97 -30 -93
rect -12 -97 -10 -93
rect -2 -97 0 -93
rect 8 -97 10 -93
rect 18 -97 20 -93
rect -22 -105 -20 -101
rect 38 -97 40 -93
rect 28 -105 30 -101
rect 78 -99 80 -93
rect 88 -97 90 -93
rect 68 -108 70 -104
rect 108 -101 110 -93
rect 118 -101 120 -93
<< ptransistor >>
rect -22 -71 -20 -65
rect -62 -81 -60 -75
rect -52 -81 -50 -75
rect -42 -81 -40 -75
rect -32 -81 -30 -75
rect 28 -71 30 -65
rect -12 -81 -10 -75
rect -2 -81 0 -75
rect 8 -81 10 -75
rect 18 -81 20 -75
rect 38 -81 40 -75
rect 68 -70 70 -64
rect 78 -81 80 -75
rect 88 -81 90 -75
rect 108 -81 110 -69
rect 118 -81 120 -69
<< ndiffusion >>
rect -63 -97 -62 -93
rect -60 -97 -59 -93
rect -53 -97 -52 -93
rect -50 -97 -49 -93
rect -43 -97 -42 -93
rect -40 -97 -39 -93
rect -33 -97 -32 -93
rect -30 -97 -29 -93
rect -13 -97 -12 -93
rect -10 -97 -9 -93
rect -3 -97 -2 -93
rect 0 -97 1 -93
rect 7 -97 8 -93
rect 10 -97 11 -93
rect 17 -97 18 -93
rect 20 -97 21 -93
rect -19 -101 -14 -97
rect -27 -105 -22 -101
rect -20 -105 -14 -101
rect -27 -109 -23 -105
rect 37 -97 38 -93
rect 40 -97 47 -93
rect 23 -105 28 -101
rect 30 -105 31 -101
rect 23 -109 27 -105
rect 41 -102 47 -97
rect 71 -95 78 -93
rect 71 -99 72 -95
rect 77 -99 78 -95
rect 80 -97 82 -93
rect 87 -97 88 -93
rect 90 -97 91 -93
rect 80 -99 84 -97
rect 66 -105 68 -104
rect 61 -108 68 -105
rect 70 -108 76 -104
rect 71 -112 76 -108
rect 107 -101 108 -93
rect 110 -101 111 -93
rect 117 -101 118 -93
rect 120 -101 121 -93
<< pdiffusion >>
rect -23 -71 -22 -65
rect -20 -71 -14 -65
rect -63 -81 -62 -75
rect -60 -81 -59 -75
rect -53 -81 -52 -75
rect -50 -81 -49 -75
rect -43 -81 -42 -75
rect -40 -81 -39 -75
rect -33 -81 -32 -75
rect -30 -81 -29 -75
rect -19 -75 -14 -71
rect 27 -71 28 -65
rect 30 -70 31 -65
rect 30 -71 37 -70
rect -13 -81 -12 -75
rect -10 -81 -9 -75
rect -3 -81 -2 -75
rect 0 -81 1 -75
rect 7 -81 8 -75
rect 10 -81 11 -75
rect 17 -81 18 -75
rect 20 -81 21 -75
rect 41 -75 47 -72
rect 37 -81 38 -75
rect 40 -81 47 -75
rect 71 -64 76 -60
rect 67 -70 68 -64
rect 70 -70 76 -64
rect 71 -80 73 -75
rect 77 -80 78 -75
rect 71 -81 78 -80
rect 80 -81 82 -75
rect 87 -81 88 -75
rect 90 -81 91 -75
rect 107 -81 108 -69
rect 110 -81 111 -69
rect 117 -81 118 -69
rect 120 -81 121 -69
<< ndcontact >>
rect -69 -97 -63 -93
rect -59 -97 -53 -93
rect -49 -97 -43 -93
rect -39 -97 -33 -93
rect -29 -97 -23 -93
rect -19 -97 -13 -93
rect -9 -97 -3 -93
rect 1 -97 7 -93
rect 11 -97 17 -93
rect 21 -97 26 -93
rect 31 -97 37 -93
rect 41 -107 47 -102
rect -27 -113 -23 -109
rect 23 -113 27 -109
rect 61 -105 66 -101
rect 72 -99 77 -95
rect 82 -97 87 -93
rect 101 -101 107 -93
rect 121 -101 127 -93
rect 71 -116 76 -112
<< pdcontact >>
rect 71 -60 77 -56
rect -29 -71 -23 -65
rect -69 -81 -63 -75
rect -59 -81 -53 -75
rect -49 -81 -43 -75
rect -39 -81 -33 -75
rect -29 -81 -23 -75
rect 21 -71 27 -65
rect -19 -81 -13 -75
rect -9 -81 -3 -75
rect 1 -81 7 -75
rect 11 -81 17 -75
rect 21 -81 26 -75
rect 41 -72 47 -67
rect 31 -81 37 -75
rect 61 -70 67 -64
rect 73 -80 77 -75
rect 82 -81 87 -75
rect 101 -81 107 -69
rect 121 -81 127 -69
<< psubstratepcontact >>
rect -10 -118 8 -112
rect 43 -118 61 -112
rect 97 -118 115 -112
<< nsubstratencontact >>
rect -10 -61 8 -55
rect 43 -60 61 -54
rect 97 -60 115 -54
<< polysilicon >>
rect -72 -109 -70 -63
rect -62 -65 -60 -63
rect -52 -65 -50 -63
rect -62 -75 -60 -71
rect -52 -75 -50 -71
rect -42 -75 -40 -63
rect -32 -75 -30 -63
rect -22 -65 -20 -62
rect -12 -65 -10 -63
rect -2 -65 0 -63
rect -62 -84 -60 -81
rect -52 -84 -50 -81
rect -42 -84 -40 -81
rect -62 -93 -60 -90
rect -52 -93 -50 -90
rect -42 -93 -40 -90
rect -32 -93 -30 -81
rect -22 -84 -20 -71
rect -12 -75 -10 -71
rect -2 -75 0 -71
rect 8 -75 10 -63
rect 18 -75 20 -63
rect 28 -65 30 -62
rect -12 -84 -10 -81
rect -2 -84 0 -81
rect 8 -84 10 -81
rect -62 -101 -60 -97
rect -52 -101 -50 -97
rect -62 -109 -60 -107
rect -52 -109 -50 -107
rect -42 -109 -40 -97
rect -32 -100 -30 -97
rect -22 -101 -20 -90
rect -12 -93 -10 -90
rect -2 -93 0 -90
rect 8 -93 10 -90
rect 18 -93 20 -81
rect 28 -84 30 -71
rect 38 -75 40 -63
rect 38 -84 40 -81
rect -12 -101 -10 -97
rect -2 -101 0 -97
rect -32 -109 -30 -105
rect -22 -109 -20 -105
rect -12 -109 -10 -107
rect -2 -108 0 -107
rect 8 -108 10 -97
rect 18 -100 20 -97
rect 28 -101 30 -90
rect 38 -93 40 -90
rect 18 -108 20 -105
rect 28 -108 30 -105
rect 38 -108 40 -97
rect 48 -110 50 -63
rect 58 -110 60 -62
rect 68 -64 70 -61
rect 78 -67 80 -62
rect 88 -66 90 -62
rect 68 -80 70 -70
rect 78 -75 80 -72
rect 88 -75 90 -71
rect 78 -84 80 -81
rect 88 -84 90 -81
rect 68 -104 70 -84
rect 78 -93 80 -90
rect 88 -93 90 -90
rect 78 -102 80 -99
rect 88 -103 90 -97
rect 68 -111 70 -108
rect 78 -110 80 -107
rect 88 -110 90 -108
rect 98 -110 100 -62
rect 108 -69 110 -62
rect 118 -69 120 -62
rect 108 -84 110 -81
rect 118 -84 120 -81
rect 108 -93 110 -90
rect 118 -93 120 -90
rect 108 -110 110 -101
rect 118 -110 120 -101
rect 128 -110 130 -62
<< polycontact >>
rect -42 -90 -38 -84
rect -24 -90 -20 -84
rect 8 -90 12 -84
rect 28 -90 32 -84
rect 66 -84 70 -80
rect 106 -90 112 -84
rect 116 -90 122 -84
<< metal1 >>
rect -76 -54 134 -52
rect -76 -55 43 -54
rect -76 -60 -10 -55
rect -39 -75 -33 -60
rect -29 -65 -23 -60
rect 8 -60 43 -55
rect 61 -56 97 -54
rect 61 -60 71 -56
rect 77 -60 97 -56
rect 115 -60 134 -54
rect 11 -75 17 -60
rect 21 -65 27 -60
rect 41 -67 47 -60
rect 56 -70 61 -64
rect 67 -70 68 -64
rect -69 -83 -63 -81
rect -69 -93 -63 -91
rect -59 -88 -53 -81
rect -50 -81 -49 -75
rect -50 -93 -45 -81
rect -29 -84 -23 -81
rect -38 -90 -24 -84
rect -29 -93 -23 -90
rect -17 -93 -13 -81
rect -50 -97 -49 -93
rect -40 -97 -39 -93
rect -9 -86 -3 -81
rect -9 -93 -3 -91
rect 0 -81 1 -75
rect 29 -81 31 -75
rect 37 -80 41 -75
rect 37 -81 47 -80
rect 0 -93 5 -81
rect 21 -84 25 -81
rect 29 -84 33 -81
rect 12 -90 18 -84
rect 32 -90 33 -84
rect 21 -93 25 -90
rect 29 -93 33 -90
rect 0 -97 1 -93
rect 10 -97 11 -93
rect 29 -97 31 -93
rect 37 -94 47 -93
rect 37 -97 41 -94
rect -40 -112 -36 -97
rect -76 -113 -27 -112
rect 10 -112 14 -97
rect 29 -98 41 -97
rect 56 -94 62 -70
rect 101 -69 107 -60
rect 121 -69 127 -60
rect 77 -80 79 -75
rect 61 -99 62 -94
rect 77 -99 79 -95
rect 82 -84 87 -81
rect 82 -90 106 -84
rect 112 -90 116 -84
rect 82 -93 87 -90
rect 56 -101 62 -99
rect 56 -105 61 -101
rect -23 -113 -10 -112
rect -76 -118 -10 -113
rect 8 -113 23 -112
rect 41 -112 47 -107
rect 101 -112 107 -101
rect 121 -112 127 -101
rect 27 -113 43 -112
rect 8 -118 43 -113
rect 61 -116 71 -112
rect 76 -116 97 -112
rect 61 -118 97 -116
rect 115 -118 134 -112
rect -76 -120 134 -118
<< pm12contact >>
rect -63 -71 -58 -65
rect -54 -71 -49 -65
rect -13 -71 -8 -65
rect -4 -71 1 -65
rect 36 -90 42 -84
rect -63 -107 -58 -101
rect -54 -107 -49 -101
rect -33 -105 -28 -100
rect -13 -107 -8 -101
rect -4 -107 1 -101
rect 77 -72 82 -67
rect 86 -71 91 -66
rect 17 -105 22 -100
rect 77 -107 82 -102
rect 86 -108 91 -103
<< pdm12contact >>
rect 31 -70 37 -65
rect 91 -81 97 -75
rect 111 -81 117 -69
<< ndm12contact >>
rect 91 -99 97 -93
rect 111 -101 117 -93
rect 31 -106 37 -101
<< metal2 >>
rect -64 -61 37 -55
rect -64 -65 -58 -61
rect -4 -65 2 -61
rect -64 -71 -63 -65
rect 1 -71 2 -65
rect 7 -65 37 -61
rect -33 -100 -28 -98
rect -49 -107 -48 -101
rect -54 -111 -48 -107
rect -14 -107 -13 -101
rect -14 -111 -8 -107
rect 7 -111 13 -65
rect 56 -71 77 -66
rect 27 -80 36 -74
rect 30 -90 36 -80
rect 56 -94 61 -71
rect 74 -72 77 -71
rect 17 -100 22 -99
rect 31 -111 37 -106
rect 65 -102 70 -80
rect 91 -93 97 -81
rect 65 -107 77 -102
rect -63 -117 37 -111
<< m3contact >>
rect -49 -71 -43 -65
rect -19 -71 -13 -65
rect -33 -98 -28 -93
rect -69 -107 -63 -101
rect -4 -101 2 -96
rect 19 -80 27 -72
rect 91 -71 96 -66
rect 17 -99 22 -94
rect 111 -93 121 -81
rect 91 -108 96 -103
<< m123contact >>
rect -69 -91 -63 -83
rect -59 -93 -53 -88
rect -9 -91 -3 -86
rect 41 -80 47 -75
rect 18 -90 25 -84
rect 41 -99 47 -94
rect 56 -99 61 -94
rect 65 -80 70 -75
rect 74 -95 79 -80
<< metal3 >>
rect -49 -61 47 -55
rect -49 -65 -43 -61
rect -19 -65 -13 -61
rect 41 -75 47 -61
rect 65 -71 91 -66
rect 65 -75 70 -71
rect -9 -86 14 -83
rect -3 -88 14 -86
rect -59 -97 -33 -93
rect 9 -94 14 -88
rect 25 -90 74 -84
rect 9 -98 17 -94
rect 11 -99 17 -98
rect -4 -103 2 -101
rect 41 -103 47 -99
rect -63 -107 47 -103
rect -69 -109 47 -107
rect 56 -103 61 -99
rect 56 -108 91 -103
<< labels >>
rlabel m123contact -6 -88 -6 -88 1 transm23_out
rlabel metal1 -56 -86 -56 -86 1 transm01_out
rlabel pdm12contact 34 -68 34 -68 1 _clk
rlabel m3contact 23 -73 23 -73 1 clk
rlabel metal1 -71 -56 -71 -56 4 Vdd
rlabel metal1 -72 -115 -72 -115 2 Gnd
rlabel metal1 31 -92 31 -92 1 _nclk
rlabel metal3 48 -87 48 -87 1 nq
rlabel m123contact -66 -87 -66 -87 1 d
rlabel metal1 84 -88 84 -88 1 mux_out
rlabel metal1 82 -116 82 -116 1 Gnd
rlabel metal1 118 -56 118 -56 7 Vdd
rlabel m123contact 67 -78 67 -78 1 enable
rlabel m3contact 115 -88 115 -88 1 Q
rlabel m123contact 76 -87 76 -87 1 in_1
rlabel metal2 94 -86 94 -86 1 in_0
<< end >>
