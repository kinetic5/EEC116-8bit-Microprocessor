magic
tech scmos
timestamp 1575613539
<< nwell >>
rect 9 41 243 78
<< ntransistor >>
rect 20 29 22 35
rect 30 29 32 35
rect 40 29 42 35
rect 60 31 62 35
rect 70 29 72 35
rect 80 29 82 35
rect 100 29 102 35
rect 110 29 112 35
rect 120 29 122 35
rect 140 31 142 35
rect 150 29 152 35
rect 160 29 162 35
rect 180 26 182 35
rect 190 29 192 35
rect 200 29 202 35
rect 220 26 222 35
rect 230 26 232 35
<< ptransistor >>
rect 20 47 22 56
rect 30 47 32 56
rect 40 47 42 56
rect 60 47 62 53
rect 70 47 72 56
rect 80 47 82 56
rect 100 47 102 56
rect 110 47 112 56
rect 120 47 122 56
rect 140 47 142 53
rect 150 47 152 56
rect 160 47 162 56
rect 180 47 182 59
rect 190 47 192 56
rect 200 47 202 56
rect 220 50 222 62
rect 230 50 232 62
<< ndiffusion >>
rect 19 29 20 35
rect 22 29 23 35
rect 29 29 30 35
rect 32 30 33 35
rect 39 30 40 35
rect 32 29 40 30
rect 42 29 43 35
rect 53 34 60 35
rect 59 31 60 34
rect 62 34 70 35
rect 62 31 63 34
rect 69 29 70 34
rect 72 29 80 35
rect 82 29 83 35
rect 99 29 100 35
rect 102 29 103 35
rect 109 29 110 35
rect 112 30 113 35
rect 119 30 120 35
rect 112 29 120 30
rect 122 29 123 35
rect 133 34 140 35
rect 139 31 140 34
rect 142 34 150 35
rect 142 31 143 34
rect 149 29 150 34
rect 152 29 160 35
rect 162 29 163 35
rect 179 26 180 35
rect 182 26 183 35
rect 189 29 190 35
rect 192 29 200 35
rect 202 29 203 35
rect 219 26 220 35
rect 222 26 230 35
rect 232 28 233 35
rect 232 26 239 28
<< pdiffusion >>
rect 19 47 20 56
rect 22 47 23 56
rect 29 47 30 56
rect 32 55 40 56
rect 32 47 33 55
rect 39 47 40 55
rect 42 47 43 56
rect 59 48 60 53
rect 53 47 60 48
rect 62 51 63 53
rect 69 51 70 56
rect 62 47 70 51
rect 72 48 73 56
rect 79 48 80 56
rect 72 47 80 48
rect 82 47 83 56
rect 99 47 100 56
rect 102 47 103 56
rect 109 47 110 56
rect 112 55 120 56
rect 112 47 113 55
rect 119 47 120 55
rect 122 47 123 56
rect 139 48 140 53
rect 133 47 140 48
rect 142 51 143 53
rect 149 51 150 56
rect 142 47 150 51
rect 152 48 153 56
rect 159 48 160 56
rect 152 47 160 48
rect 162 47 163 56
rect 173 56 180 59
rect 179 47 180 56
rect 182 56 186 59
rect 182 47 183 56
rect 189 47 190 56
rect 192 47 193 56
rect 199 47 200 56
rect 202 47 203 56
rect 216 59 220 62
rect 219 50 220 59
rect 222 60 230 62
rect 222 50 223 60
rect 229 50 230 60
rect 232 59 236 62
rect 232 50 233 59
<< ndcontact >>
rect 14 29 19 35
rect 23 29 29 35
rect 43 29 49 35
rect 53 30 59 34
rect 63 29 69 34
rect 83 29 89 35
rect 93 29 99 35
rect 103 29 109 35
rect 123 29 129 35
rect 133 30 139 34
rect 143 29 149 34
rect 163 29 169 35
rect 173 26 179 35
rect 183 26 189 35
rect 203 29 209 35
rect 213 26 219 35
rect 233 28 239 35
<< pdcontact >>
rect 15 47 19 56
rect 23 47 29 56
rect 43 47 49 56
rect 63 51 69 56
rect 83 47 89 56
rect 93 47 99 56
rect 103 47 109 56
rect 123 47 129 56
rect 143 51 149 56
rect 163 47 169 56
rect 173 47 179 56
rect 183 47 189 56
rect 193 47 199 56
rect 203 47 209 56
rect 213 50 219 59
rect 223 50 229 60
rect 233 50 237 59
<< polysilicon >>
rect 10 20 12 66
rect 20 56 22 66
rect 30 65 32 66
rect 40 65 42 66
rect 30 56 32 59
rect 40 56 42 59
rect 20 44 22 47
rect 30 44 32 47
rect 40 44 42 47
rect 20 35 22 38
rect 30 35 32 38
rect 40 35 42 38
rect 20 20 22 29
rect 30 26 32 29
rect 40 26 42 29
rect 30 20 32 21
rect 40 20 42 21
rect 50 20 52 66
rect 60 53 62 66
rect 70 56 72 66
rect 80 56 82 66
rect 60 43 62 47
rect 70 43 72 47
rect 80 44 82 47
rect 60 35 62 37
rect 70 35 72 37
rect 80 35 82 38
rect 60 20 62 31
rect 70 20 72 29
rect 80 20 82 29
rect 90 20 92 66
rect 100 56 102 66
rect 110 65 112 66
rect 120 65 122 66
rect 110 56 112 59
rect 120 56 122 59
rect 100 44 102 47
rect 110 44 112 47
rect 120 44 122 47
rect 100 35 102 39
rect 110 35 112 38
rect 120 35 122 38
rect 100 20 102 29
rect 110 26 112 29
rect 120 26 122 29
rect 110 20 112 21
rect 120 20 122 21
rect 130 20 132 66
rect 140 53 142 66
rect 150 56 152 66
rect 160 56 162 66
rect 140 43 142 47
rect 150 43 152 47
rect 160 44 162 47
rect 140 35 142 37
rect 150 35 152 37
rect 160 35 162 38
rect 140 20 142 31
rect 150 20 152 29
rect 160 20 162 29
rect 170 20 172 66
rect 180 59 182 66
rect 190 56 192 59
rect 200 56 202 66
rect 180 44 182 47
rect 180 35 182 38
rect 190 35 192 47
rect 200 35 202 47
rect 180 20 182 26
rect 190 20 192 29
rect 200 26 202 29
rect 200 20 202 21
rect 210 20 212 66
rect 220 62 222 66
rect 230 62 232 66
rect 220 46 222 50
rect 230 46 232 50
rect 220 35 222 39
rect 230 35 232 39
rect 220 20 222 26
rect 230 20 232 26
rect 240 20 242 66
<< polycontact >>
rect 39 21 44 26
rect 60 37 64 43
rect 68 37 72 43
rect 119 21 124 26
rect 140 37 144 43
rect 148 37 152 43
rect 189 59 194 66
rect 180 38 184 44
<< metal1 >>
rect 6 70 208 78
rect 216 70 246 78
rect 14 56 19 70
rect 63 56 69 70
rect 83 56 89 70
rect 29 47 30 56
rect 26 35 30 47
rect 43 46 49 47
rect 43 35 49 40
rect 29 29 30 35
rect 52 48 53 53
rect 52 34 57 48
rect 93 56 99 70
rect 143 56 149 70
rect 163 56 169 70
rect 180 59 186 70
rect 182 56 186 59
rect 203 56 209 70
rect 109 47 110 56
rect 64 37 68 43
rect 106 35 110 47
rect 123 46 129 47
rect 123 35 129 40
rect 52 30 53 34
rect 14 18 19 29
rect 52 26 57 30
rect 44 21 57 26
rect 63 18 69 29
rect 109 29 110 35
rect 132 48 133 53
rect 132 34 137 48
rect 172 47 173 56
rect 182 47 183 56
rect 213 59 219 70
rect 233 59 238 70
rect 172 44 177 47
rect 193 44 199 47
rect 144 37 148 43
rect 164 38 177 44
rect 184 38 209 44
rect 172 35 177 38
rect 203 35 209 38
rect 132 30 133 34
rect 93 18 99 29
rect 132 26 137 30
rect 124 21 137 26
rect 143 18 149 29
rect 172 26 173 35
rect 183 18 189 26
rect 213 18 219 26
rect 6 10 208 18
rect 216 10 246 18
<< m2contact >>
rect 63 43 69 48
rect 83 23 89 29
rect 143 43 149 48
rect 223 60 229 67
rect 163 23 169 29
rect 233 22 239 28
<< pm12contact >>
rect 28 59 34 65
rect 38 59 44 65
rect 18 38 23 44
rect 108 59 114 65
rect 118 59 124 65
rect 78 38 83 44
rect 98 39 103 44
rect 29 21 34 26
rect 158 38 164 44
rect 218 39 223 46
rect 228 39 233 46
rect 108 21 114 26
rect 198 21 204 26
<< pdm12contact >>
rect 33 47 39 55
rect 53 48 59 55
rect 73 48 79 56
rect 113 47 119 55
rect 133 48 139 55
rect 153 48 159 56
<< ndm12contact >>
rect 33 30 39 35
rect 113 30 119 35
<< metal2 >>
rect 8 26 14 72
rect 63 66 69 80
rect 38 65 69 66
rect 44 60 69 65
rect 87 62 93 70
rect 192 70 200 78
rect 118 65 149 66
rect 63 48 69 60
rect 73 56 93 62
rect 124 60 149 65
rect 33 35 39 47
rect 53 43 63 44
rect 53 38 69 43
rect 53 26 59 38
rect 87 29 93 56
rect 143 48 149 60
rect 153 56 177 62
rect 113 35 119 47
rect 133 43 143 44
rect 89 23 93 29
rect 98 30 113 35
rect 133 38 149 43
rect 153 38 158 44
rect 171 39 177 56
rect 181 52 187 70
rect 229 60 243 67
rect 237 46 243 60
rect 98 19 104 30
rect 133 26 139 38
rect 153 34 159 38
rect 171 29 177 33
rect 169 23 177 29
rect 237 28 243 40
rect 239 21 243 28
rect 63 13 104 19
rect 63 8 69 13
rect 224 10 232 18
<< m3contact >>
rect 6 72 14 80
rect 22 59 28 65
rect 87 70 93 76
rect 181 70 187 76
rect 43 50 53 55
rect 102 59 108 65
rect 23 38 29 44
rect 73 38 78 44
rect 39 30 45 36
rect 123 50 133 55
rect 103 39 109 45
rect 8 20 15 26
rect 34 20 40 26
rect 53 20 59 26
rect 181 46 187 52
rect 218 46 224 52
rect 114 20 120 26
rect 133 20 139 26
rect 171 33 177 39
rect 227 33 233 39
rect 237 40 243 46
rect 204 22 212 29
<< m123contact >>
rect 208 70 216 78
rect 43 40 49 46
rect 123 40 129 46
rect 194 59 200 66
rect 153 23 159 34
rect 208 10 216 18
<< metal3 >>
rect 93 70 181 76
rect 200 70 208 78
rect 22 56 28 59
rect 102 56 108 59
rect 22 55 53 56
rect 22 50 43 55
rect 102 55 133 56
rect 102 50 123 55
rect 187 46 218 52
rect 6 44 43 46
rect 6 40 23 44
rect 29 40 43 44
rect 49 44 78 46
rect 49 40 73 44
rect 103 45 123 46
rect 109 40 123 45
rect 129 40 159 46
rect 243 40 246 46
rect 45 30 69 36
rect 63 26 69 30
rect 153 34 159 40
rect 15 20 25 26
rect 40 20 53 26
rect 63 20 114 26
rect 120 20 133 26
rect 177 33 227 39
rect 163 23 204 29
rect 19 16 25 20
rect 163 16 169 23
rect 212 23 243 29
rect 6 8 14 14
rect 19 10 169 16
rect 216 10 224 18
rect 237 14 243 23
rect 237 8 246 14
<< m4contact >>
rect 192 70 200 78
rect 224 10 232 18
<< m345contact >>
rect 200 59 207 66
<< metal5 >>
rect 6 59 200 66
rect 207 59 246 66
<< m456contact >>
rect 200 70 208 78
rect 216 10 224 18
<< labels >>
rlabel metal2 67 78 67 78 5 p
rlabel metal2 36 38 36 38 1 xor0_out
rlabel metal2 66 9 66 9 1 z
rlabel m3contact 241 43 241 43 7 cout
rlabel metal3 16 43 16 43 1 cin
rlabel m345contact 203 63 203 63 1 y
rlabel metal1 240 74 240 74 7 Vdd
rlabel m3contact 13 23 13 23 1 x
<< end >>
