magic
tech scmos
timestamp 1575779281
<< ntransistor >>
rect 30 30 32 34
rect 40 30 42 34
rect 60 28 62 34
rect 70 25 72 34
rect 80 28 82 34
rect 90 28 92 34
rect 110 28 112 34
rect 130 28 132 34
rect 140 28 142 34
rect 160 25 162 34
<< ptransistor >>
rect 30 46 32 52
rect 40 46 42 52
rect 60 46 62 55
rect 70 46 72 58
rect 80 46 82 55
rect 90 46 92 55
rect 110 46 112 55
rect 130 46 132 52
rect 140 46 142 52
rect 160 46 162 58
<< ndiffusion >>
rect 29 30 30 34
rect 32 30 40 34
rect 42 33 49 34
rect 42 30 43 33
rect 53 33 60 34
rect 59 28 60 33
rect 62 28 63 34
rect 69 25 70 34
rect 72 28 73 34
rect 79 28 80 34
rect 82 29 83 34
rect 89 29 90 34
rect 82 28 90 29
rect 92 28 93 34
rect 72 25 76 28
rect 109 28 110 34
rect 112 28 113 34
rect 129 28 130 34
rect 132 28 140 34
rect 142 33 149 34
rect 142 28 143 33
rect 159 25 160 34
rect 162 25 163 34
<< pdiffusion >>
rect 29 46 30 52
rect 32 47 33 52
rect 39 47 40 52
rect 32 46 40 47
rect 42 46 43 52
rect 59 47 60 55
rect 53 46 60 47
rect 62 46 63 55
rect 69 46 70 58
rect 72 55 76 58
rect 72 46 73 55
rect 79 46 80 55
rect 82 52 90 55
rect 82 46 83 52
rect 89 46 90 52
rect 92 52 96 55
rect 92 46 93 52
rect 103 54 110 55
rect 109 46 110 54
rect 112 46 113 55
rect 129 46 130 52
rect 132 47 133 52
rect 139 47 140 52
rect 132 46 140 47
rect 142 46 143 52
rect 159 46 160 58
rect 162 46 163 58
<< ndcontact >>
rect 23 28 29 34
rect 63 25 69 34
rect 73 28 79 34
rect 93 28 99 34
rect 103 28 109 34
rect 113 28 119 34
rect 123 28 129 34
rect 153 25 159 34
rect 163 25 169 34
<< pdcontact >>
rect 23 46 29 52
rect 43 46 49 52
rect 63 46 69 58
rect 73 46 79 55
rect 93 46 99 52
rect 113 46 119 55
rect 123 46 129 52
rect 143 46 149 52
rect 153 46 159 58
rect 163 46 169 58
<< polysilicon >>
rect 20 19 22 67
rect 30 52 32 67
rect 40 52 42 67
rect 30 43 32 46
rect 40 43 42 46
rect 30 34 32 37
rect 40 34 42 37
rect 30 19 32 28
rect 40 19 42 28
rect 50 19 52 67
rect 60 55 62 67
rect 70 58 72 67
rect 80 63 82 67
rect 90 63 92 67
rect 60 43 62 46
rect 70 43 72 46
rect 80 43 82 46
rect 90 43 92 46
rect 60 34 62 37
rect 70 34 72 37
rect 80 34 82 37
rect 90 34 92 37
rect 60 19 62 28
rect 70 19 72 25
rect 80 19 82 20
rect 90 19 92 20
rect 100 19 102 67
rect 110 63 112 67
rect 110 55 112 58
rect 110 43 112 46
rect 110 34 112 37
rect 110 19 112 28
rect 120 19 122 67
rect 130 52 132 67
rect 140 52 142 67
rect 130 43 132 46
rect 140 43 142 46
rect 130 34 132 37
rect 140 34 142 37
rect 130 19 132 28
rect 140 19 142 28
rect 150 19 152 67
rect 160 58 162 67
rect 160 43 162 46
rect 160 34 162 37
rect 160 19 162 25
rect 170 19 172 67
rect 180 19 182 67
rect 190 19 192 67
rect 200 19 202 67
rect 210 19 212 67
rect 220 19 222 67
rect 230 19 232 67
rect 240 19 242 67
<< polycontact >>
rect 28 37 34 43
rect 88 58 94 63
rect 58 37 63 43
rect 88 20 94 25
rect 108 58 114 63
rect 110 37 114 43
rect 128 37 134 43
<< polypplus >>
rect 80 55 82 58
rect 90 55 92 58
<< polynplus >>
rect 30 28 32 30
rect 40 28 42 30
rect 80 25 82 28
rect 90 25 92 28
<< metal1 >>
rect 6 69 208 77
rect 216 69 246 77
rect 23 52 29 69
rect 43 52 49 69
rect 63 58 69 69
rect 94 58 108 63
rect 123 55 129 69
rect 79 46 80 55
rect 23 37 28 43
rect 76 34 80 46
rect 93 34 99 40
rect 23 17 29 28
rect 79 28 80 34
rect 102 46 103 54
rect 119 52 129 55
rect 119 46 123 52
rect 143 52 149 69
rect 153 58 159 69
rect 169 46 174 58
rect 102 34 107 46
rect 167 45 174 46
rect 120 37 128 43
rect 167 39 169 45
rect 167 34 174 39
rect 102 28 103 34
rect 119 28 123 34
rect 102 25 109 28
rect 63 17 69 25
rect 94 20 109 25
rect 123 17 129 28
rect 169 25 174 34
rect 153 17 159 25
rect 6 9 208 17
rect 216 9 246 17
<< m2contact >>
rect 114 58 120 64
rect 17 37 23 43
rect 114 37 120 43
<< pm12contact >>
rect 78 58 84 63
rect 38 37 44 43
rect 68 37 73 43
rect 138 37 144 43
rect 158 37 164 43
rect 78 20 84 25
<< pdm12contact >>
rect 33 47 39 53
rect 53 47 59 55
rect 83 46 89 52
rect 103 46 109 54
rect 133 47 139 53
<< ndm12contact >>
rect 43 27 49 33
rect 53 27 59 33
rect 83 29 89 34
rect 143 27 149 33
<< metal2 >>
rect 14 71 23 77
rect 17 43 23 71
rect 63 73 69 79
rect 63 67 120 73
rect 192 69 200 77
rect 114 64 120 67
rect 43 58 49 59
rect 17 26 23 37
rect 27 33 33 53
rect 84 58 109 62
rect 78 56 109 58
rect 43 43 49 52
rect 103 54 109 56
rect 59 47 68 53
rect 44 37 49 43
rect 62 33 68 47
rect 27 27 37 33
rect 59 27 68 33
rect 83 35 89 46
rect 114 43 120 58
rect 83 34 94 35
rect 89 29 94 34
rect 88 16 94 29
rect 114 26 120 37
rect 63 10 94 16
rect 63 7 69 10
rect 224 9 232 17
<< m3contact >>
rect 6 71 14 79
rect 43 52 49 58
rect 73 37 79 43
rect 37 27 43 33
rect 127 47 133 53
rect 132 37 138 43
rect 153 37 158 43
rect 17 20 23 26
rect 72 20 78 26
rect 149 27 155 33
rect 114 20 120 26
<< m123contact >>
rect 208 69 216 77
rect 53 37 58 43
rect 93 40 99 46
rect 169 39 180 45
rect 208 9 216 17
<< metal3 >>
rect 200 69 208 77
rect 133 47 155 53
rect 37 37 53 43
rect 79 40 93 43
rect 149 43 155 47
rect 99 40 132 43
rect 79 37 132 40
rect 149 37 153 43
rect 180 39 246 45
rect 37 33 43 37
rect 149 33 155 37
rect 23 20 41 23
rect 78 20 114 26
rect 197 22 243 28
rect 17 17 41 20
rect 35 15 41 17
rect 197 15 203 22
rect 6 7 14 13
rect 35 9 203 15
rect 216 9 224 17
rect 237 13 243 22
rect 237 7 246 13
<< m4contact >>
rect 192 69 200 77
rect 224 9 232 17
<< m345contact >>
rect 42 58 49 65
<< metal5 >>
rect 6 58 42 65
rect 49 58 246 65
<< m456contact >>
rect 200 69 208 77
rect 216 9 224 17
<< labels >>
rlabel metal2 66 8 66 8 1 z
rlabel m456contact 220 13 220 13 1 Gnd
rlabel metal1 240 73 240 73 7 Vdd
rlabel metal2 66 78 66 78 5 p
rlabel m3contact 10 75 10 75 3 x
rlabel metal3 244 42 244 42 7 cout
rlabel metal5 17 62 17 62 3 y
<< end >>
