magic
tech scmos
timestamp 1575960884
<< error_p >>
rect 107 668 114 669
rect 111 614 114 666
rect -5 54 -3 57
rect -2 -1 0 54
rect -2 -3 55 -1
<< metal1 >>
rect -3 666 671 668
rect -3 614 56 666
rect 111 614 223 666
rect 279 614 391 666
rect 447 614 559 666
rect 615 614 671 666
rect -3 567 671 614
rect -3 510 -2 567
rect 55 562 671 567
rect 55 510 615 562
rect 669 510 671 562
rect -3 406 671 510
rect -3 396 615 406
rect -3 339 -2 396
rect 55 354 615 396
rect 669 354 671 406
rect 55 339 671 354
rect -3 250 671 339
rect -3 225 615 250
rect -3 168 -2 225
rect 55 198 615 225
rect 669 198 671 250
rect 55 168 671 198
rect -3 111 671 168
rect -3 -3 -2 111
rect 55 94 671 111
rect 55 42 615 94
rect 669 42 671 94
rect 55 -3 671 42
rect -3 -4 671 -3
<< metal2 >>
rect -3 666 671 668
rect -3 614 56 666
rect 111 614 223 666
rect 279 614 391 666
rect 447 614 559 666
rect 615 614 671 666
rect -3 567 671 614
rect -3 510 -2 567
rect 55 562 671 567
rect 55 510 615 562
rect 669 510 671 562
rect -3 406 671 510
rect -3 396 615 406
rect -3 339 -2 396
rect 55 354 615 396
rect 669 354 671 406
rect 55 339 671 354
rect -3 250 671 339
rect -3 225 615 250
rect -3 168 -2 225
rect 55 198 615 225
rect 669 198 671 250
rect 55 168 671 198
rect -3 111 671 168
rect -3 -3 -2 111
rect 55 94 671 111
rect 55 42 615 94
rect 669 42 671 94
rect 55 -3 671 42
rect -3 -4 671 -3
<< m123contact >>
rect 56 614 110 666
rect 223 614 279 666
rect 391 614 447 666
rect 559 614 615 666
rect -2 510 55 567
rect 615 510 669 562
rect -2 339 55 396
rect 615 354 669 406
rect -2 168 55 225
rect 615 198 669 250
rect -2 54 55 111
rect 615 42 669 94
<< metal3 >>
rect -3 666 671 668
rect -3 624 56 666
rect -3 510 -2 624
rect 55 614 56 624
rect 167 614 223 666
rect 335 614 391 666
rect 503 614 559 666
rect 669 614 671 666
rect 55 562 671 614
rect 55 510 615 562
rect -3 458 615 510
rect 669 458 671 562
rect -3 453 671 458
rect -3 339 -2 453
rect 55 406 671 453
rect 55 339 615 406
rect -3 302 615 339
rect 669 302 671 406
rect -3 282 671 302
rect -3 168 -2 282
rect 55 250 671 282
rect 55 168 615 250
rect -3 147 615 168
rect 669 147 671 250
rect -3 111 671 147
rect -3 -3 -2 111
rect 55 94 671 111
rect 55 42 615 94
rect 669 42 671 94
rect 55 -3 671 42
rect -3 -4 671 -3
<< metal4 >>
rect -3 667 671 668
rect -3 625 -2 667
rect 55 666 671 667
rect 55 625 111 666
rect -3 624 111 625
rect -3 567 -2 624
rect 55 614 111 624
rect 167 614 168 666
rect 223 614 279 666
rect 391 614 447 666
rect 559 614 615 666
rect 55 567 615 614
rect -3 562 615 567
rect 669 562 671 666
rect -3 510 671 562
rect -3 396 -2 510
rect 55 406 615 510
rect 669 406 671 510
rect 55 396 671 406
rect -3 354 671 396
rect -3 339 615 354
rect -3 225 -2 339
rect 55 250 615 339
rect 669 250 671 354
rect 55 225 671 250
rect -3 198 671 225
rect -3 168 615 198
rect -3 54 -2 168
rect 55 147 615 168
rect 669 147 671 198
rect 55 146 671 147
rect 55 94 615 146
rect 669 94 671 146
rect 55 54 671 94
rect -3 -4 671 54
<< m345contact >>
rect -2 567 55 624
rect 111 614 167 666
rect 279 614 335 666
rect 447 614 503 666
rect 615 614 669 666
rect -2 396 55 453
rect 615 458 669 510
rect -2 225 55 282
rect 615 302 669 354
rect 615 147 669 198
rect -2 54 55 111
<< metal5 >>
rect -3 667 671 668
rect -3 625 -2 667
rect 55 666 671 667
rect 55 625 111 666
rect -3 624 111 625
rect -3 567 -2 624
rect 55 614 111 624
rect 167 614 168 666
rect 223 614 279 666
rect 391 614 447 666
rect 559 614 615 666
rect 55 567 615 614
rect -3 562 615 567
rect 669 562 671 666
rect -3 510 671 562
rect -3 396 -2 510
rect 55 406 615 510
rect 669 406 671 510
rect 55 396 671 406
rect -3 354 671 396
rect -3 339 615 354
rect -3 225 -2 339
rect 55 250 615 339
rect 669 250 671 354
rect 55 225 671 250
rect -3 198 671 225
rect -3 168 615 198
rect -3 54 -2 168
rect 55 147 615 168
rect 669 147 671 198
rect 55 146 671 147
rect 55 94 615 146
rect 669 94 671 146
rect 55 54 671 94
rect -3 -4 671 54
<< m456contact >>
rect -2 625 55 667
rect 168 614 223 666
rect 335 614 391 666
rect 503 614 559 666
rect 615 562 669 614
rect -2 453 55 510
rect 615 406 669 458
rect -2 282 55 339
rect 615 250 669 302
rect -2 111 55 168
rect 615 94 669 146
<< metal6 >>
rect -3 667 671 668
rect -3 625 -2 667
rect 55 666 671 667
rect 55 625 168 666
rect -3 614 168 625
rect 223 614 335 666
rect 391 614 503 666
rect 559 614 671 666
rect -3 562 615 614
rect 669 562 671 614
rect -3 510 671 562
rect -3 453 -2 510
rect 55 458 671 510
rect 55 453 615 458
rect -3 406 615 453
rect 669 406 671 458
rect -3 339 671 406
rect -3 282 -2 339
rect 55 302 671 339
rect 55 282 615 302
rect -3 250 615 282
rect 669 250 671 302
rect -3 168 671 250
rect -3 111 -2 168
rect 55 146 671 168
rect 55 111 615 146
rect -3 94 615 111
rect 669 94 671 146
rect -3 -4 671 94
<< glass >>
rect 56 56 612 612
<< end >>
