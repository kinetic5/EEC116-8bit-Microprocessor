magic
tech scmos
timestamp 1575532930
<< nwell >>
rect -43 36 195 72
<< pwell >>
rect -43 4 195 36
<< ntransistor >>
rect -30 26 -28 30
rect -20 26 -18 30
rect 0 26 2 30
rect 10 26 12 30
rect 30 26 32 30
rect 40 26 42 30
rect 60 26 62 30
rect 70 26 72 30
rect 90 26 92 30
rect 100 26 102 30
rect 120 26 122 30
rect 130 26 132 30
rect 140 26 142 30
rect 160 24 162 30
rect 170 26 172 30
rect 180 26 182 30
rect 150 16 152 22
<< ptransistor >>
rect -30 42 -28 48
rect -20 42 -18 48
rect 0 42 2 48
rect 10 42 12 48
rect 30 42 32 48
rect 40 42 42 48
rect 60 42 62 48
rect 70 42 72 48
rect 90 42 92 48
rect 100 42 102 48
rect 120 42 122 48
rect 130 42 132 48
rect 140 42 142 48
rect 150 42 152 51
rect 160 42 162 51
rect 170 42 172 48
rect 180 42 182 48
<< ndiffusion >>
rect -31 26 -30 30
rect -28 26 -20 30
rect -18 26 -17 30
rect -1 26 0 30
rect 2 26 3 30
rect 9 26 10 30
rect 12 26 13 30
rect 29 26 30 30
rect 32 26 33 30
rect 39 26 40 30
rect 42 26 43 30
rect 59 26 60 30
rect 62 26 63 30
rect 69 26 70 30
rect 72 26 73 30
rect 89 26 90 30
rect 92 26 93 30
rect 99 26 100 30
rect 102 26 103 30
rect 119 26 120 30
rect 122 26 123 30
rect 129 26 130 30
rect 132 26 140 30
rect 142 26 143 30
rect 153 24 160 30
rect 162 26 163 30
rect 169 26 170 30
rect 172 26 180 30
rect 182 26 183 30
rect 162 24 166 26
rect 153 22 159 24
rect 149 16 150 22
rect 152 16 159 22
<< pdiffusion >>
rect -37 46 -30 48
rect -31 42 -30 46
rect -28 46 -20 48
rect -28 42 -27 46
rect -21 42 -20 46
rect -18 42 -17 48
rect -1 42 0 48
rect 2 46 10 48
rect 2 42 3 46
rect 9 42 10 46
rect 12 46 16 48
rect 12 42 13 46
rect 26 46 30 48
rect 29 42 30 46
rect 32 46 40 48
rect 32 42 33 46
rect 39 42 40 46
rect 42 46 46 48
rect 42 42 43 46
rect 56 47 60 48
rect 59 42 60 47
rect 62 46 70 48
rect 62 42 63 46
rect 69 42 70 46
rect 72 46 76 48
rect 72 42 73 46
rect 86 46 90 48
rect 89 42 90 46
rect 92 46 100 48
rect 92 42 93 46
rect 99 42 100 46
rect 102 46 106 48
rect 102 42 103 46
rect 146 48 150 51
rect 116 47 120 48
rect 119 42 120 47
rect 122 46 130 48
rect 122 42 123 46
rect 129 42 130 46
rect 132 47 140 48
rect 132 42 133 47
rect 139 42 140 47
rect 142 47 150 48
rect 142 42 143 47
rect 149 42 150 47
rect 152 48 160 51
rect 152 42 153 48
rect 159 42 160 48
rect 162 48 166 51
rect 162 42 163 48
rect 169 42 170 48
rect 172 46 180 48
rect 172 42 173 46
rect 179 42 180 46
rect 182 46 189 48
rect 182 42 183 46
<< ndcontact >>
rect -37 26 -31 30
rect -17 26 -11 30
rect 3 26 9 30
rect 13 26 19 30
rect 23 26 29 30
rect 33 26 39 30
rect 43 26 48 30
rect 53 26 59 30
rect 63 26 69 30
rect 73 26 79 30
rect 83 26 89 30
rect 93 26 99 30
rect 103 26 108 30
rect 113 26 119 30
rect 123 26 129 30
rect 143 26 149 30
rect 163 26 169 30
rect 183 26 189 30
<< pdcontact >>
rect -37 42 -31 46
rect -27 42 -21 46
rect -17 42 -11 48
rect 3 42 9 46
rect 13 42 19 46
rect 23 42 29 46
rect 33 42 39 46
rect 43 42 48 46
rect 63 42 69 46
rect 73 42 79 46
rect 83 42 89 46
rect 93 42 99 46
rect 103 42 108 46
rect 123 42 129 46
rect 133 42 139 47
rect 143 42 149 47
rect 163 42 169 48
rect 173 42 179 46
rect 183 42 189 46
<< psubstratepcontact >>
rect -36 13 -31 18
rect 1 7 6 12
rect 32 7 37 12
rect 59 7 64 12
rect 85 7 90 12
rect 111 7 116 12
rect 138 7 143 12
rect 163 7 168 12
rect 187 7 192 12
<< nsubstratencontact >>
rect -31 64 -26 69
rect 0 64 5 69
rect 30 64 35 69
rect 55 64 60 69
rect 91 64 96 69
rect 116 64 121 69
rect 175 64 180 69
rect 164 59 169 64
<< polysilicon >>
rect -40 15 -38 54
rect -30 48 -28 50
rect -20 48 -18 54
rect -30 30 -28 42
rect -20 30 -18 42
rect -30 15 -28 26
rect -20 23 -18 26
rect -20 15 -18 16
rect -10 15 -8 54
rect 0 48 2 54
rect 10 48 12 54
rect 0 39 2 42
rect 10 39 12 42
rect 0 30 2 33
rect 10 30 12 34
rect 0 15 2 26
rect 10 15 12 26
rect 20 15 22 54
rect 30 48 32 49
rect 40 48 42 50
rect 30 39 32 42
rect 40 39 42 42
rect 30 30 32 33
rect 40 30 42 33
rect 30 23 32 26
rect 40 23 42 26
rect 30 15 32 18
rect 40 15 42 19
rect 50 15 52 53
rect 60 48 62 50
rect 70 48 72 54
rect 60 38 62 42
rect 70 39 72 42
rect 60 30 62 33
rect 70 30 72 34
rect 60 15 62 26
rect 70 15 72 26
rect 80 15 82 54
rect 90 48 92 49
rect 100 48 102 50
rect 90 39 92 42
rect 100 39 102 42
rect 90 30 92 33
rect 100 30 102 33
rect 90 23 92 26
rect 100 23 102 26
rect 90 15 92 18
rect 100 13 102 19
rect 110 13 112 54
rect 120 48 122 50
rect 130 48 132 54
rect 150 51 152 54
rect 160 51 162 54
rect 140 48 142 50
rect 170 48 172 54
rect 180 48 182 49
rect 120 38 122 42
rect 120 30 122 33
rect 130 30 132 42
rect 140 30 142 42
rect 150 38 152 42
rect 120 13 122 26
rect 130 23 132 26
rect 130 13 132 18
rect 140 13 142 26
rect 150 22 152 32
rect 160 39 162 42
rect 160 30 162 33
rect 170 30 172 42
rect 180 30 182 42
rect 150 13 152 16
rect 160 13 162 24
rect 170 21 172 26
rect 180 13 182 26
rect 190 13 192 54
<< polycontact >>
rect -30 50 -26 54
rect -2 33 3 39
rect 40 50 44 54
rect 40 19 44 23
rect 58 50 62 54
rect 100 50 104 54
rect 100 19 104 23
rect 118 50 122 54
rect 147 32 152 38
rect 160 33 165 39
<< metal1 >>
rect -40 69 133 72
rect -40 64 -31 69
rect -26 64 0 69
rect 5 64 30 69
rect 35 64 55 69
rect 60 64 91 69
rect 96 64 116 69
rect 121 64 133 69
rect 141 64 149 72
rect 157 64 165 72
rect 173 69 192 72
rect 173 64 175 69
rect 180 64 192 69
rect -37 46 -33 64
rect -26 50 -22 54
rect -17 48 -11 64
rect 3 46 9 64
rect 40 54 62 55
rect 44 51 58 54
rect 19 42 23 46
rect -27 39 -21 42
rect -27 33 -2 39
rect -17 30 -11 33
rect 23 30 29 42
rect -37 18 -31 26
rect 19 26 23 30
rect 33 36 39 42
rect 33 31 34 36
rect 33 30 39 31
rect 43 39 48 42
rect 43 30 48 34
rect 52 42 54 47
rect 65 46 70 64
rect 104 51 118 54
rect 69 42 70 46
rect 79 42 83 46
rect 52 30 56 42
rect 83 30 89 42
rect 52 26 53 30
rect 69 26 70 30
rect 79 26 83 30
rect 93 36 99 42
rect 93 31 94 36
rect 93 30 99 31
rect 103 39 108 42
rect 103 30 108 34
rect 112 42 114 47
rect 125 46 130 64
rect 145 47 149 64
rect 163 59 164 64
rect 163 48 169 59
rect 129 42 130 46
rect 185 46 189 64
rect 112 30 116 42
rect 133 38 139 42
rect 173 39 179 42
rect 133 33 147 38
rect 143 32 147 33
rect 165 33 189 39
rect 143 30 149 32
rect 183 30 189 33
rect 112 26 113 30
rect 122 26 123 30
rect -37 13 -36 18
rect -37 12 -31 13
rect 3 12 9 26
rect 52 23 56 26
rect 44 19 56 23
rect 65 12 70 26
rect 112 23 116 26
rect 104 19 116 23
rect 122 12 127 26
rect 163 12 167 26
rect -40 4 -28 12
rect -20 4 -12 12
rect -4 7 1 12
rect 6 7 32 12
rect 37 7 59 12
rect 64 7 85 12
rect 90 7 111 12
rect 116 7 138 12
rect 143 7 163 12
rect 168 7 187 12
rect -4 4 192 7
<< m2contact >>
rect 43 34 48 39
rect 103 34 108 39
<< pm12contact >>
rect 30 49 35 54
rect 9 34 14 39
rect 90 49 95 54
rect 59 33 64 38
rect 69 34 74 39
rect 137 50 142 55
rect 177 49 182 54
rect 119 33 124 38
rect -24 16 -18 23
rect 29 18 34 23
rect 89 18 94 23
rect 130 18 135 23
rect 170 15 176 21
<< pdm12contact >>
rect -7 42 -1 48
rect 54 42 59 47
rect 114 42 119 47
rect 153 42 159 48
<< ndm12contact >>
rect -7 24 -1 30
rect 143 16 149 22
<< metal2 >>
rect -36 23 -31 67
rect -18 48 -13 67
rect 54 47 59 49
rect -7 39 -1 42
rect -7 30 -1 34
rect 9 39 14 40
rect 69 45 74 74
rect 114 47 119 49
rect 43 39 48 40
rect 9 19 14 34
rect 69 39 74 40
rect 103 39 108 40
rect 20 14 25 31
rect 29 23 34 27
rect 124 33 129 67
rect 133 50 137 55
rect 133 45 138 50
rect 119 28 135 33
rect 119 27 124 28
rect 89 23 94 27
rect 130 23 135 28
rect 153 22 159 42
rect 177 36 182 49
rect 149 16 159 22
rect 20 9 74 14
rect 69 2 74 9
<< m3contact >>
rect -36 67 -31 72
rect -18 67 -13 72
rect 35 49 40 54
rect 54 49 59 54
rect -20 42 -13 48
rect -7 34 -1 39
rect 9 40 14 45
rect 43 40 48 45
rect 124 67 129 72
rect 95 49 100 54
rect 114 49 119 54
rect -36 18 -31 23
rect -18 16 -12 23
rect 20 31 25 36
rect 69 40 74 45
rect 103 40 108 45
rect 9 13 15 19
rect 34 22 39 27
rect 59 22 64 33
rect 133 40 138 45
rect 159 42 165 48
rect 94 22 99 27
rect 119 22 124 27
rect 177 31 182 36
rect 164 15 170 21
<< m123contact >>
rect -27 54 -22 59
rect 34 31 39 36
rect 94 31 99 36
rect 133 64 141 72
rect 149 64 157 72
rect 165 64 173 72
rect -28 4 -20 12
rect -12 4 -4 12
<< metal3 >>
rect -40 67 -36 72
rect -13 67 124 72
rect 185 67 192 74
rect -40 59 128 63
rect -40 58 -27 59
rect -22 58 128 59
rect 123 57 128 58
rect 183 58 192 63
rect 183 57 188 58
rect 40 49 54 54
rect 100 49 114 54
rect 123 52 188 57
rect -40 42 -20 48
rect 14 40 43 45
rect 74 40 103 45
rect 108 40 133 45
rect 165 42 192 48
rect 9 39 14 40
rect -1 34 14 39
rect 25 31 34 36
rect 59 33 94 36
rect -31 18 -18 23
rect -12 18 5 23
rect 39 22 59 27
rect 64 31 94 33
rect 99 31 133 36
rect 128 30 133 31
rect 177 30 182 31
rect 99 22 119 27
rect 128 25 182 30
rect 0 9 5 18
rect 15 15 164 18
rect 15 13 170 15
rect 0 4 192 9
rect 185 2 192 4
<< m4contact >>
rect 141 64 149 72
rect 157 64 165 72
rect -36 4 -28 12
rect -20 4 -12 12
<< metal4 >>
rect 149 64 157 72
rect -28 4 -20 12
<< labels >>
rlabel metal2 72 73 72 73 5 p
rlabel metal2 22 10 22 10 1 z
rlabel ndm12contact 146 19 146 19 1 cout
rlabel metal3 11 36 11 36 1 and_gate_to_xor_nand
rlabel metal3 61 36 61 36 1 xor1_to_xor2_nand
rlabel metal1 145 37 145 37 1 p_cin_nand_to_nand_cout
rlabel metal3 -39 60 -39 60 3 y
rlabel metal3 -9 70 -9 70 5 cin
rlabel metal4 153 68 153 68 1 Vdd
rlabel metal4 -24 8 -24 8 1 Gnd
rlabel m3contact -34 71 -34 71 4 x
<< end >>
