magic
tech scmos
timestamp 1575939707
<< metal1 >>
rect 0 0 667 667
<< metal2 >>
rect 0 0 667 667
<< metal3 >>
rect 0 0 667 667
<< metal4 >>
rect 0 0 667 667
<< metal5 >>
rect 0 0 667 667
<< metal6 >>
rect 0 0 667 667
<< end >>
