magic
tech scmos
timestamp 1575939553
<< metal1 >>
rect 247 70 487 78
rect 474 18 480 19
rect 247 10 487 18
<< ndm12contact >>
rect 284 25 290 31
<< metal2 >>
rect 284 18 290 25
rect 284 17 291 18
rect 284 11 310 17
rect 304 8 310 11
<< metal3 >>
rect 269 38 300 47
rect 275 37 300 38
rect 275 36 293 37
rect 285 17 293 36
rect 247 8 255 14
rect 285 11 487 17
rect 478 8 487 11
<< metal5 >>
rect 247 59 497 66
use and  and_0
timestamp 1575855885
transform 1 0 251 0 1 6
box 0 4 42 72
use inputff  inputff_0
timestamp 1575939406
transform -1 0 421 0 1 130
box -76 -120 134 -52
<< labels >>
rlabel metal5 253 62 253 62 1 y
rlabel metal2 307 9 307 9 1 z
rlabel metal1 485 74 485 74 7 Vdd
<< end >>
