magic
tech scmos
timestamp 1575427599
<< ntransistor >>
rect -30 28 -28 32
rect -20 28 -18 32
rect 0 28 2 32
rect 10 28 12 32
rect 30 28 32 32
rect 40 28 42 32
rect 60 28 62 32
rect 70 28 72 32
rect 90 28 92 32
rect 100 28 102 32
rect 120 28 122 32
rect 130 28 132 32
rect 140 28 142 32
rect 160 28 162 32
rect 170 28 172 32
rect 180 28 182 32
rect 150 20 152 24
<< ptransistor >>
rect -30 44 -28 50
rect -20 44 -18 50
rect 0 44 2 50
rect 10 44 12 50
rect 30 44 32 50
rect 40 44 42 50
rect 60 44 62 50
rect 70 44 72 50
rect 90 44 92 50
rect 100 44 102 50
rect 120 44 122 50
rect 130 44 132 50
rect 140 44 142 50
rect 150 44 152 50
rect 160 44 162 50
rect 170 44 172 50
rect 180 44 182 50
<< ndiffusion >>
rect -31 28 -30 32
rect -28 28 -20 32
rect -18 28 -17 32
rect -1 28 0 32
rect 2 28 3 32
rect 9 28 10 32
rect 12 28 13 32
rect 29 28 30 32
rect 32 28 33 32
rect 39 28 40 32
rect 42 28 43 32
rect 59 28 60 32
rect 62 28 63 32
rect 69 28 70 32
rect 72 28 73 32
rect 89 28 90 32
rect 92 28 93 32
rect 99 28 100 32
rect 102 28 103 32
rect 119 28 120 32
rect 122 28 123 32
rect 129 28 130 32
rect 132 28 140 32
rect 142 28 143 32
rect 154 28 160 32
rect 162 28 163 32
rect 169 28 170 32
rect 172 28 180 32
rect 182 28 183 32
rect 154 24 158 28
rect 149 20 150 24
rect 152 20 158 24
<< pdiffusion >>
rect -37 48 -30 50
rect -31 44 -30 48
rect -28 48 -20 50
rect -28 44 -27 48
rect -21 44 -20 48
rect -18 44 -17 50
rect -1 44 0 50
rect 2 48 10 50
rect 2 44 3 48
rect 9 44 10 48
rect 12 48 16 50
rect 12 44 13 48
rect 26 48 30 50
rect 29 44 30 48
rect 32 48 40 50
rect 32 44 33 48
rect 39 44 40 48
rect 42 48 46 50
rect 42 44 43 48
rect 56 49 60 50
rect 59 44 60 49
rect 62 48 70 50
rect 62 44 63 48
rect 69 44 70 48
rect 72 48 76 50
rect 72 44 73 48
rect 86 48 90 50
rect 89 44 90 48
rect 92 48 100 50
rect 92 44 93 48
rect 99 44 100 48
rect 102 48 106 50
rect 102 44 103 48
rect 116 49 120 50
rect 119 44 120 49
rect 122 48 130 50
rect 122 44 123 48
rect 129 44 130 48
rect 132 49 140 50
rect 132 44 133 49
rect 139 44 140 49
rect 142 49 150 50
rect 142 44 143 49
rect 149 44 150 49
rect 152 44 153 50
rect 159 44 160 50
rect 162 48 170 50
rect 162 44 163 48
rect 169 44 170 48
rect 172 48 180 50
rect 172 44 173 48
rect 179 44 180 48
rect 182 48 189 50
rect 182 44 183 48
<< ndcontact >>
rect -37 28 -31 32
rect -17 28 -11 32
rect 3 28 9 32
rect 13 28 19 32
rect 23 28 29 32
rect 33 28 39 32
rect 43 28 48 32
rect 53 28 59 32
rect 63 28 69 32
rect 73 28 79 32
rect 83 28 89 32
rect 93 28 99 32
rect 103 28 108 32
rect 113 28 119 32
rect 123 28 129 32
rect 143 28 149 32
rect 163 28 169 32
rect 183 28 189 32
<< pdcontact >>
rect -37 44 -31 48
rect -27 44 -21 48
rect -17 44 -11 50
rect 3 44 9 48
rect 13 44 19 48
rect 23 44 29 48
rect 33 44 39 48
rect 43 44 48 48
rect 63 44 69 48
rect 73 44 79 48
rect 83 44 89 48
rect 93 44 99 48
rect 103 44 108 48
rect 123 44 129 48
rect 133 44 139 49
rect 143 44 149 49
rect 163 44 169 48
rect 173 44 179 48
rect 183 44 189 48
<< polysilicon >>
rect -40 17 -38 56
rect -30 50 -28 52
rect -20 50 -18 56
rect -30 32 -28 44
rect -20 32 -18 44
rect -30 17 -28 28
rect -20 25 -18 28
rect -10 17 -8 56
rect 0 50 2 56
rect 10 50 12 56
rect 0 41 2 44
rect 10 41 12 44
rect 0 32 2 35
rect 10 32 12 36
rect 0 17 2 28
rect 10 17 12 28
rect 20 17 22 56
rect 30 50 32 51
rect 40 50 42 52
rect 30 41 32 44
rect 40 41 42 44
rect 30 32 32 35
rect 40 32 42 35
rect 30 25 32 28
rect 40 25 42 28
rect 30 17 32 20
rect 40 17 42 21
rect 50 17 52 55
rect 60 50 62 52
rect 70 50 72 56
rect 60 40 62 44
rect 70 41 72 44
rect 60 32 62 35
rect 70 32 72 36
rect 60 17 62 28
rect 70 17 72 28
rect 80 17 82 56
rect 90 50 92 51
rect 100 50 102 52
rect 90 41 92 44
rect 100 41 102 44
rect 90 32 92 35
rect 100 32 102 35
rect 90 25 92 28
rect 100 25 102 28
rect 90 17 92 20
rect 100 17 102 21
rect 110 17 112 56
rect 120 50 122 52
rect 130 50 132 56
rect 140 50 142 52
rect 150 50 152 56
rect 160 50 162 56
rect 170 50 172 56
rect 180 50 182 51
rect 120 40 122 44
rect 120 32 122 35
rect 130 32 132 44
rect 140 32 142 44
rect 150 41 152 44
rect 120 17 122 28
rect 130 25 132 28
rect 130 17 132 20
rect 140 17 142 28
rect 150 24 152 34
rect 160 41 162 44
rect 160 32 162 35
rect 170 32 172 44
rect 180 32 182 44
rect 150 17 152 20
rect 160 17 162 28
rect 170 23 172 28
rect 180 17 182 28
rect 190 17 192 56
<< polycontact >>
rect -30 52 -26 56
rect -2 35 3 41
rect 40 52 44 56
rect 40 21 44 25
rect 58 52 62 56
rect 100 52 104 56
rect 100 21 104 25
rect 118 52 122 56
rect 147 34 152 41
rect 160 35 165 41
<< metal1 >>
rect -40 66 192 74
rect -37 48 -33 66
rect -17 50 -11 66
rect 3 48 9 66
rect 40 56 62 57
rect 44 53 58 56
rect 19 44 23 48
rect -27 41 -21 44
rect -27 35 -2 41
rect -17 32 -11 35
rect 23 32 29 44
rect -37 10 -31 28
rect 19 28 23 32
rect 33 38 39 44
rect 33 33 34 38
rect 33 32 39 33
rect 43 41 48 44
rect 43 32 48 36
rect 52 44 54 49
rect 65 48 70 66
rect 104 53 118 56
rect 69 44 70 48
rect 79 44 83 48
rect 52 32 56 44
rect 83 32 89 44
rect 52 28 53 32
rect 69 28 70 32
rect 79 28 83 32
rect 93 38 99 44
rect 93 33 94 38
rect 93 32 99 33
rect 103 41 108 44
rect 103 32 108 36
rect 112 44 114 49
rect 125 48 130 66
rect 145 49 149 66
rect 129 44 130 48
rect 163 48 169 66
rect 185 48 189 66
rect 112 32 116 44
rect 133 41 139 44
rect 173 41 179 44
rect 133 35 147 41
rect 143 34 147 35
rect 165 35 189 41
rect 143 32 149 34
rect 183 32 189 35
rect 112 28 113 32
rect 122 28 123 32
rect 3 10 9 28
rect 52 25 56 28
rect 44 21 56 25
rect 65 10 70 28
rect 112 25 116 28
rect 104 21 116 25
rect 122 10 127 28
rect 163 10 167 28
rect -40 2 192 10
<< m2contact >>
rect 43 36 48 41
rect 103 36 108 41
<< pm12contact >>
rect 30 51 35 56
rect 9 36 14 41
rect 90 51 95 56
rect 59 35 64 40
rect 69 36 74 41
rect 137 52 142 57
rect 177 51 182 56
rect 119 35 124 40
rect -24 17 -18 25
rect 29 20 34 25
rect 89 20 94 25
rect 130 20 135 25
rect 170 17 176 23
<< pdm12contact >>
rect -7 44 -1 50
rect 54 44 59 49
rect 114 44 119 49
rect 153 44 159 50
<< ndm12contact >>
rect -7 26 -1 32
rect 143 18 149 24
<< metal2 >>
rect -40 9 -35 69
rect -20 50 -13 69
rect -20 43 -13 44
rect 54 49 59 51
rect -7 41 -1 44
rect -7 32 -1 36
rect 9 41 14 42
rect 69 47 74 76
rect 114 49 119 51
rect 43 41 48 42
rect 9 17 14 36
rect 69 41 74 42
rect 103 41 108 42
rect 20 16 25 33
rect 124 35 129 69
rect 133 52 137 57
rect 133 47 138 52
rect 59 25 64 30
rect 119 30 135 35
rect 119 25 124 30
rect 130 25 135 30
rect 153 24 159 44
rect 177 38 182 51
rect 149 18 159 24
rect 20 11 74 16
rect 69 0 74 11
<< m3contact >>
rect -40 69 -33 76
rect -20 69 -13 74
rect 35 51 40 56
rect 54 51 59 56
rect -20 44 -13 50
rect -7 36 -1 41
rect 9 42 14 47
rect 43 42 48 47
rect 124 69 129 74
rect 95 51 100 56
rect 114 51 119 56
rect -24 11 -18 17
rect 20 33 25 38
rect 69 42 74 47
rect 103 42 108 47
rect 9 11 15 17
rect 59 30 64 35
rect 133 42 138 47
rect 153 50 159 56
rect 34 20 39 25
rect 59 20 64 25
rect 94 20 99 25
rect 119 20 124 25
rect 177 33 182 38
rect 170 11 176 17
rect -40 2 -33 9
<< m123contact >>
rect -30 56 -24 63
rect 34 33 39 38
rect 94 33 99 38
<< metal3 >>
rect -13 69 124 74
rect 185 69 192 76
rect -40 63 192 65
rect -40 60 -30 63
rect -24 60 192 63
rect 40 51 54 56
rect 100 51 114 56
rect -40 44 -20 50
rect 14 42 43 47
rect 74 42 103 47
rect 108 42 133 47
rect 153 44 192 50
rect 9 41 14 42
rect -1 36 14 41
rect 25 33 34 38
rect 59 35 94 38
rect 64 33 94 35
rect 99 33 177 38
rect 39 20 59 25
rect 99 20 119 25
rect 15 11 170 16
rect -24 7 -18 11
rect -33 2 192 7
<< labels >>
rlabel metal1 3 6 3 6 2 Gnd
rlabel metal2 22 12 22 12 1 z
rlabel ndm12contact 146 21 146 21 1 cout
rlabel metal3 -9 72 -9 72 5 cin
rlabel metal2 72 75 72 75 5 p
rlabel metal3 -39 62 -39 62 3 y
rlabel m3contact -38 71 -38 71 4 x
rlabel metal3 11 38 11 38 1 and_gate_to_xor_nand
rlabel metal3 61 38 61 38 1 xor1_to_xor2_nand
rlabel metal1 145 39 145 39 1 p_cin_nand_to_nand_cout
rlabel metal1 -28 70 -28 70 1 Vdd
<< end >>
