magic
tech scmos
timestamp 1575690611
<< nwell >>
rect -52 -20 154 16
<< pwell >>
rect -52 -56 154 -20
<< ntransistor >>
rect -40 -35 -38 -31
rect -30 -35 -28 -31
rect -10 -35 -8 -31
rect 0 -35 2 -31
rect 20 -35 22 -31
rect 30 -35 32 -31
rect 40 -43 42 -39
rect 60 -35 62 -31
rect 70 -35 72 -31
rect 80 -35 82 -31
rect 90 -35 92 -31
rect 120 -35 122 -31
rect 130 -35 132 -31
rect 100 -43 102 -39
rect 140 -43 142 -39
<< ptransistor >>
rect -40 -11 -38 -5
rect -30 -11 -28 -5
rect -10 -11 -8 -5
rect 0 -11 2 -5
rect 40 -2 42 3
rect 20 -11 22 -5
rect 30 -11 32 -5
rect 100 -2 102 3
rect 60 -11 62 -5
rect 70 -11 72 -5
rect 80 -11 82 -5
rect 90 -11 92 -5
rect 140 -2 142 3
rect 120 -11 122 -5
rect 130 -11 132 -5
<< ndiffusion >>
rect -41 -35 -40 -31
rect -38 -35 -37 -31
rect -31 -35 -30 -31
rect -28 -35 -27 -31
rect -11 -35 -10 -31
rect -8 -35 -7 -31
rect -1 -35 0 -31
rect 2 -35 3 -31
rect 19 -35 20 -31
rect 22 -35 24 -31
rect 28 -35 30 -31
rect 32 -35 33 -31
rect 34 -43 35 -39
rect 39 -43 40 -39
rect 42 -43 45 -39
rect 54 -35 55 -31
rect 59 -35 60 -31
rect 62 -35 64 -31
rect 69 -35 70 -31
rect 72 -35 74 -31
rect 78 -35 80 -31
rect 82 -35 83 -31
rect 89 -35 90 -31
rect 92 -35 94 -31
rect 118 -35 120 -31
rect 122 -35 123 -31
rect 129 -35 130 -31
rect 132 -35 134 -31
rect 94 -43 95 -39
rect 99 -43 100 -39
rect 102 -43 104 -39
rect 139 -43 140 -39
rect 142 -43 144 -39
<< pdiffusion >>
rect -41 -11 -40 -5
rect -38 -11 -37 -5
rect -31 -11 -30 -5
rect -28 -11 -27 -5
rect -11 -11 -10 -5
rect -8 -11 -6 -5
rect -2 -11 0 -5
rect 2 -6 7 -5
rect 2 -11 3 -6
rect 34 -1 35 3
rect 39 -1 40 3
rect 34 -2 40 -1
rect 42 -2 44 3
rect 14 -6 20 -5
rect 19 -11 20 -6
rect 22 -11 24 -5
rect 28 -11 30 -5
rect 32 -6 38 -5
rect 32 -11 34 -6
rect 94 -1 95 3
rect 99 -1 100 3
rect 94 -2 100 -1
rect 102 -2 104 3
rect 54 -11 55 -5
rect 59 -11 60 -5
rect 62 -11 63 -5
rect 69 -11 70 -5
rect 72 -11 73 -5
rect 79 -11 80 -5
rect 82 -11 83 -5
rect 89 -11 90 -5
rect 92 -6 98 -5
rect 92 -11 94 -6
rect 139 -1 140 3
rect 134 -2 140 -1
rect 142 -2 144 3
rect 118 -11 120 -5
rect 122 -11 123 -5
rect 129 -11 130 -5
rect 132 -6 138 -5
rect 132 -11 134 -6
<< ndcontact >>
rect -46 -35 -41 -31
rect -37 -35 -31 -31
rect -27 -35 -22 -31
rect -15 -35 -11 -31
rect -7 -35 -1 -31
rect 3 -35 7 -31
rect 15 -35 19 -31
rect 24 -35 28 -31
rect 33 -35 37 -31
rect 35 -43 39 -39
rect 45 -43 49 -39
rect 55 -35 59 -31
rect 64 -35 69 -31
rect 74 -35 78 -31
rect 83 -35 89 -31
rect 94 -35 98 -31
rect 114 -35 118 -31
rect 123 -35 129 -31
rect 134 -35 138 -31
rect 95 -43 99 -39
rect 104 -43 108 -39
rect 134 -43 139 -39
rect 144 -43 148 -39
<< pdcontact >>
rect -46 -11 -41 -5
rect -37 -11 -31 -5
rect -27 -11 -22 -5
rect -15 -11 -11 -5
rect -6 -11 -2 -5
rect 3 -11 7 -6
rect 35 -1 39 3
rect 44 -2 48 3
rect 24 -11 28 -5
rect 34 -11 38 -6
rect 95 -1 99 3
rect 104 -2 108 3
rect 55 -11 59 -5
rect 63 -11 69 -5
rect 73 -11 79 -5
rect 83 -11 89 -5
rect 94 -11 98 -6
rect 134 -1 139 3
rect 144 -2 148 3
rect 114 -11 118 -5
rect 123 -11 129 -5
rect 134 -11 138 -6
<< psubstratepcontact >>
rect -27 -53 -15 -47
rect 50 -53 62 -47
rect 105 -53 117 -47
<< nsubstratencontact >>
rect -31 6 -19 13
rect 12 7 24 13
rect 57 6 69 13
rect 104 7 116 13
<< polysilicon >>
rect 20 3 22 6
rect 30 3 32 6
rect 40 3 42 6
rect -50 -43 -48 3
rect -40 -5 -38 3
rect -30 -5 -28 3
rect -40 -24 -38 -11
rect -30 -14 -28 -11
rect -40 -31 -38 -28
rect -30 -31 -28 -19
rect -40 -43 -38 -35
rect -30 -43 -28 -35
rect -20 -43 -18 3
rect -10 -5 -8 -2
rect 0 -5 2 -2
rect -10 -16 -8 -11
rect 0 -16 2 -11
rect -10 -31 -8 -26
rect 0 -31 2 -26
rect -10 -38 -8 -35
rect 0 -38 2 -35
rect 10 -43 12 3
rect 20 -5 22 -2
rect 30 -5 32 -2
rect 20 -16 22 -11
rect 30 -16 32 -11
rect 40 -24 42 -2
rect 20 -31 22 -28
rect 30 -31 32 -28
rect 20 -38 22 -35
rect 30 -38 32 -35
rect 40 -39 42 -29
rect 50 -43 52 6
rect 100 3 102 6
rect 60 -5 62 -1
rect 70 -5 72 -1
rect 80 -5 82 -2
rect 90 -5 92 -2
rect 60 -31 62 -11
rect 70 -23 72 -11
rect 80 -16 82 -11
rect 90 -16 92 -11
rect 100 -23 102 -2
rect 70 -31 72 -28
rect 80 -31 82 -28
rect 90 -31 92 -28
rect 60 -38 62 -35
rect 70 -43 72 -35
rect 80 -38 82 -35
rect 90 -38 92 -35
rect 100 -39 102 -28
rect 110 -39 112 6
rect 140 3 142 6
rect 120 -5 122 -1
rect 130 -5 132 -1
rect 120 -23 122 -11
rect 130 -23 132 -11
rect 140 -23 142 -2
rect 120 -31 122 -28
rect 130 -31 132 -28
rect 120 -39 122 -35
rect 130 -39 132 -35
rect 140 -39 142 -28
rect 150 -39 152 -1
rect 40 -46 42 -43
rect 100 -46 102 -43
rect 140 -46 142 -43
<< polycontact >>
rect -40 -28 -36 -24
rect 129 -28 133 -23
<< metal1 >>
rect -50 13 154 14
rect -50 6 -31 13
rect -19 7 12 13
rect 24 7 57 13
rect -19 6 57 7
rect 69 7 104 13
rect 116 7 154 13
rect 69 6 154 7
rect -37 -5 -31 6
rect 35 3 39 6
rect -48 -11 -46 -5
rect -22 -11 -20 -5
rect -48 -31 -43 -16
rect -25 -24 -20 -11
rect -36 -26 -20 -24
rect -36 -28 -26 -26
rect -21 -31 -20 -26
rect -48 -35 -46 -31
rect -22 -35 -20 -31
rect -16 -11 -15 -5
rect -16 -31 -13 -11
rect -6 -26 -2 -11
rect 2 -11 3 -6
rect -16 -35 -15 -31
rect 2 -31 5 -11
rect 15 -31 18 -11
rect 24 -24 28 -11
rect 34 -14 37 -11
rect 24 -31 28 -29
rect 34 -31 37 -19
rect 2 -35 3 -31
rect -37 -46 -31 -35
rect 48 -39 52 3
rect 63 -5 69 6
rect 95 3 99 6
rect 108 -2 109 3
rect 55 -14 59 -11
rect 55 -31 59 -19
rect 75 -31 78 -11
rect 83 -22 89 -11
rect 83 -31 89 -28
rect 92 -11 94 -6
rect 92 -12 98 -11
rect 92 -17 94 -12
rect 92 -31 95 -17
rect 92 -35 94 -31
rect 106 -32 109 -2
rect 123 -5 129 6
rect 134 3 139 6
rect 138 -11 140 -6
rect 114 -12 117 -11
rect 114 -31 117 -17
rect 136 -23 140 -11
rect 145 -15 148 -2
rect 145 -19 154 -15
rect 125 -28 129 -23
rect 136 -28 137 -23
rect 136 -31 140 -28
rect 49 -43 57 -39
rect 35 -46 39 -43
rect 65 -46 69 -35
rect 138 -35 140 -31
rect 105 -39 109 -37
rect 108 -43 109 -39
rect 95 -46 99 -43
rect 123 -46 129 -35
rect 145 -39 148 -19
rect 134 -46 139 -43
rect -50 -47 154 -46
rect -50 -53 -27 -47
rect -15 -53 50 -47
rect 62 -53 105 -47
rect 117 -53 154 -47
rect -50 -54 154 -53
<< m2contact >>
rect -48 -16 -43 -11
rect -26 -31 -21 -26
rect -6 -31 -1 -26
rect 34 -19 39 -14
rect 24 -29 29 -24
rect 7 -36 12 -31
rect 55 -19 60 -14
rect 83 -28 89 -22
rect 94 -17 99 -12
rect 112 -17 117 -12
rect 105 -37 110 -32
<< pm12contact >>
rect -12 -2 -7 3
rect -3 -2 2 3
rect 17 -2 22 3
rect 27 -2 32 3
rect -33 -19 -28 -14
rect 40 -29 45 -24
rect -12 -43 -7 -38
rect -3 -43 2 -38
rect 17 -43 22 -38
rect 27 -43 32 -38
rect 77 -2 82 3
rect 87 -2 92 3
rect 67 -28 72 -23
rect 98 -28 103 -23
rect 120 -28 125 -23
rect 137 -28 142 -23
rect 57 -43 62 -38
rect 77 -43 82 -38
rect 87 -43 92 -38
<< pdm12contact >>
rect 14 -11 19 -6
<< metal2 >>
rect -33 -14 -28 16
rect 17 8 92 10
rect 22 7 92 8
rect 87 3 92 7
rect 2 -2 3 3
rect 32 -2 72 3
rect -2 -13 3 -2
rect -13 -17 3 -13
rect 8 -11 14 -6
rect 27 -8 30 -2
rect 87 -5 91 -2
rect 24 -11 30 -8
rect 86 -8 91 -5
rect -26 -52 -21 -31
rect -13 -38 -10 -17
rect 8 -21 11 -11
rect 24 -15 28 -11
rect 86 -13 89 -8
rect -5 -24 11 -21
rect 16 -19 28 -15
rect 39 -19 55 -14
rect 76 -17 89 -13
rect 99 -17 112 -12
rect -5 -26 -1 -24
rect -13 -43 -12 -38
rect 16 -38 20 -19
rect 29 -29 40 -24
rect 57 -28 67 -25
rect 57 -29 72 -28
rect 57 -38 62 -29
rect 16 -43 17 -38
rect 76 -38 79 -17
rect 89 -28 98 -23
rect 142 -28 154 -23
rect 120 -32 124 -28
rect 110 -37 124 -32
rect 76 -43 77 -38
rect 17 -52 22 -43
rect 137 -47 142 -28
rect 41 -51 142 -47
rect -26 -55 22 -52
<< m3contact >>
rect -48 -11 -43 -5
rect 17 3 22 8
rect -17 -2 -12 3
rect 72 -2 77 3
rect -12 -48 -7 -43
rect 7 -41 12 -36
rect 32 -43 37 -38
rect 92 -43 97 -38
rect -3 -48 2 -43
rect 36 -52 41 -47
<< metal3 >>
rect -48 8 22 12
rect -48 7 17 8
rect -48 -5 -43 7
rect -12 -19 -7 3
rect -12 -22 2 -19
rect -3 -43 2 -22
rect -12 -56 -7 -48
rect -3 -56 2 -48
rect 7 -47 12 -41
rect 17 -38 22 3
rect 77 -2 82 3
rect 78 -13 82 -2
rect 78 -18 92 -13
rect 17 -43 32 -38
rect 87 -43 92 -18
rect 7 -52 36 -47
<< labels >>
rlabel metal1 -14 -22 -14 -22 3 D
rlabel metal1 149 -17 149 -17 7 Qbar
rlabel metal2 149 -26 149 -26 7 Q
rlabel metal2 -31 15 -31 15 5 clk
rlabel metal1 26 11 26 11 5 Vdd
rlabel metal1 4 -50 4 -50 1 Gnd
rlabel m3contact -10 -45 -10 -45 1 EN
rlabel m3contact 0 -45 0 -45 1 ENbar
<< end >>
