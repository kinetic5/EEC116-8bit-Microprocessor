magic
tech scmos
timestamp 1576013044
<< error_p >>
rect 15432 1541 15433 1545
rect 15436 1539 15437 1541
<< metal1 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1543 13975 1569
rect -1773 1541 15766 1543
rect -1773 1529 15098 1541
rect -1773 1232 -1767 1529
rect -754 1232 15098 1529
rect -1773 1214 15098 1232
rect -1773 226 -1444 1214
rect 15425 1214 15766 1541
rect 15437 1197 15766 1214
rect -1773 -623 -1772 226
rect -1449 -623 -1444 226
rect -1773 -654 -1444 -623
rect -1216 657 14878 986
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -1336 -1441 -665
rect -3013 -1341 -1441 -1336
rect -1773 -15993 -1444 -1341
rect -1216 -15423 -887 657
rect 232 650 561 657
rect 14873 645 14878 657
rect 15437 868 15441 1197
rect 232 456 561 457
rect -667 127 14661 456
rect -666 -14873 -337 127
rect -116 -95 213 -94
rect 577 -95 14100 -94
rect -116 -423 14100 -95
rect -116 -14336 213 -423
rect 13771 -3679 14100 -423
rect 13756 -4525 14100 -3679
rect 13756 -14333 14085 -4525
rect -116 -14341 222 -14336
rect 582 -14341 13655 -14336
rect -116 -14658 13655 -14341
rect -116 -14665 222 -14658
rect 588 -14665 13655 -14658
rect 14323 -14871 14655 127
rect 14873 -1424 15202 645
rect 232 -14873 561 -14872
rect 866 -14873 14655 -14871
rect -666 -14876 14655 -14873
rect -666 -15202 14211 -14876
rect -664 -15211 14211 -15202
rect 14645 -15200 14655 -14876
rect 14870 -3055 15202 -1424
rect 14870 -14709 15199 -3055
rect 15437 -13974 15766 868
rect 15434 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 14870 -15053 14871 -14709
rect 15437 -14766 15766 -14654
rect 14645 -15211 14649 -15200
rect 14870 -15418 15199 -15053
rect 232 -15423 561 -15420
rect -1216 -15752 14778 -15423
rect 15521 -14799 15766 -14766
rect 15521 -15983 15646 -14799
rect 15437 -15989 15646 -15983
rect 10 -15993 661 -15992
rect 15437 -15993 15768 -15989
rect -1773 -15998 8414 -15993
rect -1773 -16081 14470 -15998
rect -1773 -16210 15766 -16081
rect -1773 -16315 14469 -16210
rect -1773 -16322 10 -16315
rect 661 -16322 14469 -16315
rect 7835 -16324 14469 -16322
rect 15753 -16324 15766 -16210
rect 7835 -16327 15766 -16324
rect 10 -17229 661 -16553
<< metal2 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1546 13975 1569
rect 240 1543 15763 1546
rect -1774 1541 15763 1543
rect -1774 1538 15098 1541
rect -1774 1529 13299 1538
rect -1774 1232 -1767 1529
rect -754 1232 13299 1529
rect -1774 1217 13299 1232
rect -1774 1214 890 1217
rect -1774 1211 -1445 1214
rect -1774 255 -1767 1211
rect -1456 255 -1445 1211
rect 13971 1217 15098 1538
rect 15425 1219 15436 1541
rect 15758 1219 15763 1541
rect 15425 1217 15763 1219
rect 15434 1197 15763 1217
rect -929 981 14512 982
rect -1774 226 -1445 255
rect -1774 -623 -1772 226
rect -1449 -623 -1445 226
rect -1774 -654 -1445 -623
rect -1217 814 14512 981
rect -1217 664 12407 814
rect 13092 664 14512 814
rect -1217 660 14512 664
rect 14852 660 14878 982
rect -1217 653 14878 660
rect -1217 652 896 653
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -670 -1441 -665
rect -1835 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -1835 -1336 -1441 -1331
rect -3013 -1341 -1441 -1336
rect -1774 -15992 -1445 -1341
rect -1217 -1544 -888 652
rect 15434 868 15441 1197
rect 14884 618 15213 645
rect -1217 -2224 -1047 -1544
rect -889 -2224 -888 -1544
rect -1217 -15428 -888 -2224
rect -667 444 876 457
rect -667 129 14649 444
rect -667 -14001 -339 129
rect 467 116 14649 129
rect 1720 -95 2049 -94
rect 2520 -95 14096 -93
rect -116 -422 14096 -95
rect -116 -423 3442 -422
rect -116 -424 222 -423
rect 582 -424 3442 -423
rect -116 -13100 213 -424
rect 13767 -1532 14096 -422
rect 13932 -2213 14096 -1532
rect -116 -13787 42 -13100
rect 200 -13787 213 -13100
rect -667 -14674 -482 -14001
rect -116 -14333 213 -13787
rect 13767 -13979 14096 -2213
rect 14095 -14312 14096 -13979
rect 13767 -14333 14096 -14312
rect 14321 -636 14649 116
rect 14321 -1321 14327 -636
rect 14499 -1321 14649 -636
rect -116 -14341 222 -14333
rect 582 -14341 13267 -14333
rect -116 -14347 13267 -14341
rect -116 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -116 -14662 13267 -14484
rect 13646 -14662 13655 -14333
rect 14321 -14517 14649 -1321
rect 14884 -13082 15213 272
rect 15028 -13769 15213 -13082
rect -667 -14883 -339 -14674
rect 14321 -14850 14327 -14517
rect 14884 -14709 15213 -13769
rect 14321 -14876 14649 -14850
rect -667 -15043 13336 -14883
rect 14002 -15043 14211 -14883
rect -667 -15211 14211 -15043
rect 14645 -15211 14649 -14876
rect 15212 -15053 15213 -14709
rect 14884 -15063 15213 -15053
rect 15212 -15398 15213 -15063
rect 14884 -15418 15213 -15398
rect -1217 -15609 14338 -15428
rect -1217 -15757 886 -15609
rect 1567 -15757 14338 -15609
rect 14772 -15757 14778 -15428
rect 15212 -15757 15213 -15418
rect 15434 -13972 15763 868
rect 15434 -14674 15436 -13972
rect 15747 -13974 15763 -13972
rect 15747 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 15747 -14674 15763 -14654
rect 15434 -14694 15763 -14674
rect 15434 -14766 15766 -14694
rect 15521 -14771 15766 -14766
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -14799 15766 -14771
rect 15644 -15986 15646 -14799
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16081 14470 -15993
rect 662 -16090 15766 -16081
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16210 15766 -16204
rect 662 -16313 14469 -16210
rect -1774 -16315 14469 -16313
rect -1774 -16321 10 -16315
rect -9 -16322 10 -16321
rect 661 -16321 14469 -16315
rect 15753 -16321 15766 -16210
rect 10 -17229 661 -16553
<< m123contact >>
rect 13308 1569 13962 1943
rect -1767 1232 -754 1529
rect 15098 1212 15425 1541
rect -1772 -623 -1449 226
rect -2255 -1336 -1835 -665
rect 14878 645 15219 991
rect 15441 868 15768 1197
rect 13655 -14672 14099 -14333
rect 14211 -15222 14645 -14876
rect 14871 -15053 15212 -14709
rect 14778 -15764 15212 -15418
rect 15766 -14654 15975 -13974
rect 15434 -15983 15521 -14766
rect 15646 -15989 15768 -14799
rect 14470 -16081 15768 -15993
rect 10 -16553 661 -16315
rect 14469 -16324 15753 -16210
<< metal3 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1546 13975 1569
rect -1774 1541 15763 1546
rect -1774 1538 15098 1541
rect -1774 1529 13299 1538
rect -1774 1232 -1767 1529
rect -754 1232 13299 1529
rect -1774 1217 13299 1232
rect -1774 1211 -1445 1217
rect -1774 255 -1767 1211
rect -1456 255 -1445 1211
rect 13971 1217 15098 1538
rect 15425 1219 15436 1541
rect 15758 1219 15763 1541
rect 15425 1217 15763 1219
rect 15434 1197 15763 1217
rect -1774 226 -1445 255
rect -1774 -623 -1772 226
rect -1449 -623 -1445 226
rect -1774 -654 -1445 -623
rect -1224 982 1544 984
rect -1224 814 14512 982
rect -1224 664 12407 814
rect 13092 664 14512 814
rect -1224 660 14512 664
rect 14852 660 14878 982
rect -1224 655 14878 660
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -670 -1441 -665
rect -1835 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -1835 -1336 -1441 -1331
rect -3013 -1341 -1441 -1336
rect -1774 -15992 -1445 -1341
rect -1224 -1544 -895 655
rect 466 653 14878 655
rect 15434 868 15441 1197
rect 14884 618 15213 645
rect -667 444 1547 454
rect -667 125 14656 444
rect -1224 -2224 -1047 -1544
rect -1224 -15428 -895 -2224
rect -667 -14001 -338 125
rect 108 115 14656 125
rect -115 -101 2593 -94
rect -115 -423 14094 -101
rect -115 -13100 214 -423
rect 2416 -430 14094 -423
rect 13765 -1532 14094 -430
rect 13932 -2213 14094 -1532
rect -115 -13787 42 -13100
rect 200 -13787 214 -13100
rect -667 -14674 -482 -14001
rect -115 -14334 214 -13787
rect 13765 -13979 14094 -2213
rect 14327 -636 14656 115
rect 14499 -1321 14656 -636
rect 13765 -14333 14094 -14312
rect -115 -14347 13267 -14334
rect -115 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -115 -14663 13267 -14484
rect 13646 -14663 13655 -14334
rect 14327 -14517 14656 -1321
rect 14884 -13082 15213 272
rect 15028 -13769 15213 -13082
rect -667 -14889 -338 -14674
rect 14884 -14709 15213 -13769
rect 14327 -14876 14656 -14850
rect -667 -15043 13336 -14889
rect 14002 -15043 14211 -14889
rect -667 -15218 14211 -15043
rect 14645 -15218 14656 -14876
rect 15212 -15053 15213 -14709
rect 14884 -15063 15213 -15053
rect 15212 -15398 15213 -15063
rect 14884 -15418 15213 -15398
rect -1224 -15609 14338 -15428
rect -1224 -15757 886 -15609
rect 1567 -15757 14338 -15609
rect 14772 -15757 14778 -15428
rect 15212 -15757 15213 -15418
rect 15434 -13972 15763 868
rect 15434 -14674 15436 -13972
rect 15747 -13974 15763 -13972
rect 15747 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 15747 -14674 15763 -14654
rect 15434 -14694 15763 -14674
rect 15434 -14766 15766 -14694
rect 15521 -14771 15766 -14766
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -14799 15766 -14771
rect 15644 -15986 15646 -14799
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16081 14470 -15993
rect 662 -16090 15766 -16081
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16210 15766 -16204
rect 662 -16313 14469 -16210
rect -1774 -16315 14469 -16313
rect -1774 -16321 10 -16315
rect -9 -16322 10 -16321
rect 661 -16321 14469 -16315
rect 15753 -16321 15766 -16210
rect 10 -17229 661 -16553
<< m234contact >>
rect -1767 255 -1456 1211
rect 13299 1209 13971 1538
rect 15436 1219 15758 1541
rect 12407 664 13092 814
rect 14512 660 14852 987
rect -1816 -1331 -1462 -670
rect 14875 272 15216 618
rect -1047 -2224 -889 -1544
rect 13764 -2213 13932 -1532
rect 42 -13787 200 -13100
rect -482 -14674 -311 -14001
rect 14327 -1321 14499 -636
rect 13757 -14312 14095 -13979
rect 12441 -14484 13126 -14347
rect 13267 -14668 13646 -14333
rect 14872 -13769 15028 -13082
rect 14327 -14850 14665 -14517
rect 13336 -15043 14002 -14877
rect 14877 -15398 15212 -15063
rect 886 -15760 1567 -15609
rect 14338 -15757 14772 -15422
rect 15436 -14674 15747 -13972
rect 15529 -15986 15644 -14771
rect -7 -16313 662 -15992
rect 14468 -16204 15752 -16090
<< metal4 >>
rect 13304 1549 13975 2669
rect 1879 1539 15433 1549
rect 15529 1541 15770 1549
rect -1767 1538 15436 1539
rect -1767 1220 13299 1538
rect -1767 1211 8012 1220
rect -1456 1210 8012 1211
rect -1456 255 -1438 1210
rect 13971 1220 15436 1538
rect 13971 1218 13975 1220
rect 15433 1219 15436 1220
rect 15758 1220 15770 1541
rect 15758 1219 15762 1220
rect -1767 -629 -1438 255
rect -1217 984 2672 989
rect -1217 973 14512 984
rect -1217 823 12407 973
rect 13092 823 14512 973
rect -1217 814 14512 823
rect -1217 664 12407 814
rect 13092 664 14512 814
rect -1217 660 14512 664
rect 14852 660 15213 984
rect -1767 -654 -1441 -629
rect -3013 -670 -1441 -654
rect -3013 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -3013 -1341 -1441 -1331
rect -1767 -1356 -1441 -1341
rect -1767 -15992 -1438 -1356
rect -1217 -1544 -888 660
rect 1910 655 15213 660
rect 14884 618 15213 655
rect -1217 -1546 -1047 -1544
rect -1217 -2226 -1215 -1546
rect -1057 -2224 -1047 -1546
rect -889 -2224 -888 -1544
rect -1057 -2226 -888 -2224
rect -1217 -15415 -888 -2226
rect -667 451 2201 454
rect -667 125 14656 451
rect -667 -13991 -338 125
rect -322 122 14656 125
rect -667 -14664 -663 -13991
rect -492 -14001 -338 -13991
rect -115 -94 6919 -87
rect -115 -416 14094 -94
rect -115 -13096 214 -416
rect 2735 -423 14094 -416
rect 13765 -1530 14094 -423
rect 14327 -636 14656 122
rect 14499 -1321 14510 -636
rect 14327 -1323 14510 -1321
rect 13765 -1532 13945 -1530
rect 13932 -2213 13945 -1532
rect -115 -13778 -111 -13096
rect 28 -13100 214 -13096
rect 28 -13778 42 -13100
rect -115 -13787 42 -13778
rect 200 -13787 214 -13100
rect -492 -14664 -482 -14001
rect -667 -14674 -482 -14664
rect -115 -14334 214 -13787
rect 13765 -13979 14094 -2213
rect -115 -14347 13267 -14334
rect -115 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -115 -14532 13267 -14484
rect -115 -14663 12447 -14532
rect 13132 -14663 13267 -14532
rect 13765 -14334 14094 -14312
rect 13646 -14663 14094 -14334
rect 14327 -14517 14656 -1323
rect 14884 -13082 15213 272
rect 15028 -13761 15035 -13082
rect 15212 -13761 15213 -13082
rect 15028 -13769 15213 -13761
rect -667 -14882 -338 -14674
rect -667 -15043 13336 -14882
rect 14327 -14882 14656 -14850
rect 14002 -15043 14656 -14882
rect -667 -15064 14656 -15043
rect 14884 -15063 15213 -13769
rect -667 -15211 13341 -15064
rect 14007 -15211 14656 -15064
rect 15212 -15398 15213 -15063
rect 14884 -15415 15213 -15398
rect -1217 -15421 15213 -15415
rect -1217 -15598 886 -15421
rect 1567 -15422 15213 -15421
rect 1567 -15598 14338 -15422
rect -1217 -15609 14338 -15598
rect -1217 -15744 886 -15609
rect 1567 -15744 14338 -15609
rect 14772 -15744 15213 -15422
rect 15433 -13972 15762 1219
rect 15433 -14674 15436 -13972
rect 15747 -13974 15762 -13972
rect 15747 -14654 16673 -13974
rect 15747 -14674 15762 -14654
rect 15433 -14694 15762 -14674
rect 15433 -14771 15766 -14694
rect 15433 -15986 15529 -14771
rect 15644 -15986 15766 -14771
rect 15433 -15989 15766 -15986
rect 15433 -15992 15768 -15989
rect -1788 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16090 15766 -15993
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16313 15766 -16204
rect -1788 -16321 15766 -16313
rect -9 -16322 661 -16321
rect 10 -17229 661 -16322
<< metal5 >>
rect 12407 973 13089 2672
rect 12407 661 13089 823
rect 14325 -1320 14510 -640
rect 14657 -1320 16677 -640
rect -3000 -2224 -1215 -1549
rect -1057 -2224 -893 -1549
rect 13759 -2210 13945 -1533
rect 14102 -2210 16674 -1533
rect -3003 -13778 -111 -13096
rect 28 -13778 209 -13096
rect 14870 -13761 15035 -13086
rect 15212 -13761 16670 -13086
rect 14870 -13764 16670 -13761
rect -3003 -13787 209 -13778
rect -3009 -14664 -663 -13998
rect -492 -14664 -323 -13998
rect -3009 -14672 -323 -14664
rect 12444 -14532 13130 -14343
rect 12444 -14669 12447 -14532
rect 886 -15421 1565 -15415
rect 886 -17232 1565 -15598
rect 12444 -17227 13130 -14669
rect 13339 -15064 14003 -14871
rect 13339 -15230 13341 -15064
rect 13339 -17237 14003 -15230
<< m456contact >>
rect 12407 823 13092 973
rect 14510 -1323 14657 -636
rect -1215 -2226 -1057 -1546
rect 13945 -2213 14102 -1530
rect -111 -13778 28 -13096
rect 15035 -13761 15212 -13082
rect -663 -14664 -492 -13991
rect 12447 -14669 13132 -14532
rect 886 -15598 1567 -15421
rect 13341 -15230 14007 -15064
<< metal6 >>
rect 12407 973 13089 2672
rect 12407 661 13089 823
rect 14325 -1320 14510 -640
rect 14657 -1320 16677 -640
rect -3000 -2224 -1215 -1549
rect -1057 -2224 -893 -1549
rect 13759 -2210 13945 -1533
rect 14102 -2210 16674 -1533
rect -3003 -13778 -111 -13096
rect 28 -13778 209 -13096
rect 14870 -13761 15035 -13086
rect 15212 -13761 16670 -13086
rect 14870 -13764 16670 -13761
rect -3003 -13787 209 -13778
rect -3009 -14664 -663 -13998
rect -492 -14664 -323 -13998
rect -3009 -14672 -323 -14664
rect 12444 -14532 13130 -14343
rect 12444 -14669 12447 -14532
rect 886 -15421 1565 -15415
rect 886 -17232 1565 -15598
rect 12444 -17227 13130 -14669
rect 13339 -15064 14003 -14871
rect 13339 -15230 13341 -15064
rect 13339 -17237 14003 -15230
use pad  pad_48
timestamp 1575998002
transform 1 0 -29 0 1 2000
box -3 -4 672 668
use pad  pad_49
timestamp 1575998002
transform 1 0 860 0 1 2000
box -3 -4 672 668
use pad  pad_50
timestamp 1575998002
transform 1 0 1749 0 1 2000
box -3 -4 672 668
use pad  pad_51
timestamp 1575998002
transform 1 0 2638 0 1 2000
box -3 -4 672 668
use pad  pad_52
timestamp 1575998002
transform 1 0 3527 0 1 2000
box -3 -4 672 668
use pad  pad_53
timestamp 1575998002
transform 1 0 4416 0 1 2000
box -3 -4 672 668
use pad  pad_54
timestamp 1575998002
transform 1 0 5305 0 1 2000
box -3 -4 672 668
use pad  pad_55
timestamp 1575998002
transform 1 0 6194 0 1 2000
box -3 -4 672 668
use pad  pad_56
timestamp 1575998002
transform 1 0 7083 0 1 2000
box -3 -4 672 668
use pad  pad_57
timestamp 1575998002
transform 1 0 7972 0 1 2000
box -3 -4 672 668
use pad  pad_58
timestamp 1575998002
transform 1 0 8861 0 1 2000
box -3 -4 672 668
use pad  pad_59
timestamp 1575998002
transform 1 0 9750 0 1 2000
box -3 -4 672 668
use pad  pad_60
timestamp 1575998002
transform 1 0 10639 0 1 2000
box -3 -4 672 668
use pad  pad_61
timestamp 1575998002
transform 1 0 11528 0 1 2000
box -3 -4 672 668
use pad  pad_62
timestamp 1575998002
transform 1 0 12417 0 1 2000
box -3 -4 672 668
use pad  pad_63
timestamp 1575998002
transform 1 0 13306 0 1 2000
box -3 -4 672 668
use pad  pad_32
timestamp 1575998002
transform 0 1 -2998 -1 0 -662
box -3 -4 672 668
use pad  pad_16
timestamp 1575998002
transform 0 1 16001 -1 0 -645
box -3 -4 672 668
use pad  pad_33
timestamp 1575998002
transform 0 1 -2998 -1 0 -1551
box -3 -4 672 668
use pad  pad_17
timestamp 1575998002
transform 0 1 16001 -1 0 -1534
box -3 -4 672 668
use pad  pad_34
timestamp 1575998002
transform 0 1 -2998 -1 0 -2440
box -3 -4 672 668
use pad  pad_18
timestamp 1575998002
transform 0 1 16001 -1 0 -2423
box -3 -4 672 668
use pad  pad_35
timestamp 1575998002
transform 0 1 -2998 -1 0 -3329
box -3 -4 672 668
use pad  pad_19
timestamp 1575998002
transform 0 1 16001 -1 0 -3312
box -3 -4 672 668
use pad  pad_36
timestamp 1575998002
transform 0 1 -2998 -1 0 -4218
box -3 -4 672 668
use pad  pad_20
timestamp 1575998002
transform 0 1 16001 -1 0 -4201
box -3 -4 672 668
use pad  pad_37
timestamp 1575998002
transform 0 1 -2998 -1 0 -5107
box -3 -4 672 668
use pad  pad_21
timestamp 1575998002
transform 0 1 16001 -1 0 -5090
box -3 -4 672 668
use pad  pad_38
timestamp 1575998002
transform 0 1 -2998 -1 0 -5996
box -3 -4 672 668
use pad  pad_22
timestamp 1575998002
transform 0 1 16001 -1 0 -5979
box -3 -4 672 668
use pad  pad_39
timestamp 1575998002
transform 0 1 -2998 -1 0 -6885
box -3 -4 672 668
use pad  pad_23
timestamp 1575998002
transform 0 1 16001 -1 0 -6868
box -3 -4 672 668
use pad  pad_40
timestamp 1575998002
transform 0 1 -2998 -1 0 -7774
box -3 -4 672 668
use pad  pad_24
timestamp 1575998002
transform 0 1 16001 -1 0 -7757
box -3 -4 672 668
use pad  pad_41
timestamp 1575998002
transform 0 1 -2998 -1 0 -8663
box -3 -4 672 668
use pad  pad_25
timestamp 1575998002
transform 0 1 16001 -1 0 -8646
box -3 -4 672 668
use pad  pad_42
timestamp 1575998002
transform 0 1 -2998 -1 0 -9552
box -3 -4 672 668
use pad  pad_26
timestamp 1575998002
transform 0 1 16001 -1 0 -9535
box -3 -4 672 668
use pad  pad_43
timestamp 1575998002
transform 0 1 -2998 -1 0 -10441
box -3 -4 672 668
use pad  pad_27
timestamp 1575998002
transform 0 1 16001 -1 0 -10424
box -3 -4 672 668
use pad  pad_44
timestamp 1575998002
transform 0 1 -2998 -1 0 -11330
box -3 -4 672 668
use pad  pad_28
timestamp 1575998002
transform 0 1 16001 -1 0 -11313
box -3 -4 672 668
use pad  pad_45
timestamp 1575998002
transform 0 1 -2998 -1 0 -12219
box -3 -4 672 668
use pad  pad_29
timestamp 1575998002
transform 0 1 16001 -1 0 -12202
box -3 -4 672 668
use pad  pad_46
timestamp 1575998002
transform 0 1 -2998 -1 0 -13108
box -3 -4 672 668
use pad  pad_30
timestamp 1575998002
transform 0 1 16001 -1 0 -13091
box -3 -4 672 668
use pad  pad_47
timestamp 1575998002
transform 0 1 -2998 -1 0 -13997
box -3 -4 672 668
use pad  pad_31
timestamp 1575998002
transform 0 1 16001 -1 0 -13980
box -3 -4 672 668
use pad  pad_0
timestamp 1575998002
transform 1 0 0 0 1 -17223
box -3 -4 672 668
use pad  pad_1
timestamp 1575998002
transform 1 0 889 0 1 -17223
box -3 -4 672 668
use pad  pad_2
timestamp 1575998002
transform 1 0 1778 0 1 -17223
box -3 -4 672 668
use pad  pad_3
timestamp 1575998002
transform 1 0 2667 0 1 -17223
box -3 -4 672 668
use pad  pad_4
timestamp 1575998002
transform 1 0 3556 0 1 -17223
box -3 -4 672 668
use pad  pad_5
timestamp 1575998002
transform 1 0 4445 0 1 -17223
box -3 -4 672 668
use pad  pad_6
timestamp 1575998002
transform 1 0 5334 0 1 -17223
box -3 -4 672 668
use pad  pad_7
timestamp 1575998002
transform 1 0 6223 0 1 -17223
box -3 -4 672 668
use pad  pad_8
timestamp 1575998002
transform 1 0 7112 0 1 -17223
box -3 -4 672 668
use pad  pad_9
timestamp 1575998002
transform 1 0 8001 0 1 -17223
box -3 -4 672 668
use pad  pad_10
timestamp 1575998002
transform 1 0 8890 0 1 -17223
box -3 -4 672 668
use pad  pad_11
timestamp 1575998002
transform 1 0 9779 0 1 -17223
box -3 -4 672 668
use pad  pad_12
timestamp 1575998002
transform 1 0 10668 0 1 -17223
box -3 -4 672 668
use pad  pad_13
timestamp 1575998002
transform 1 0 11557 0 1 -17223
box -3 -4 672 668
use pad  pad_14
timestamp 1575998002
transform 1 0 12446 0 1 -17223
box -3 -4 672 668
use pad  pad_15
timestamp 1575998002
transform 1 0 13335 0 1 -17223
box -3 -4 672 668
<< labels >>
rlabel metal4 6989 -16182 6989 -16182 1 VddIo
rlabel metal4 7131 -15637 7131 -15637 1 GndIo
rlabel metal4 7143 -15058 7143 -15058 1 VddCore
rlabel metal4 7143 -14490 7143 -14490 1 GndCore
<< end >>
