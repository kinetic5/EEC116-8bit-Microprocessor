magic
tech scmos
timestamp 1575941163
<< error_p >>
rect 55 613 56 667
rect 228 613 229 667
rect 393 613 394 667
rect 558 613 559 667
rect 54 612 55 613
rect 0 605 55 606
rect 613 549 666 550
rect 0 440 55 441
rect 613 384 666 385
rect 0 275 55 276
rect 613 219 666 220
rect 0 110 55 111
rect 613 54 666 55
rect 165 1 166 54
rect 330 1 331 54
rect 495 1 496 54
rect 612 53 613 54
<< metal1 >>
rect 0 613 118 667
rect 173 613 283 667
rect 338 613 448 667
rect 503 613 613 667
rect 0 604 613 613
rect 0 550 666 604
rect 55 495 666 550
rect 0 494 666 495
rect 0 439 613 494
rect 0 385 666 439
rect 55 330 666 385
rect 0 329 666 330
rect 0 274 613 329
rect 0 220 666 274
rect 55 165 666 220
rect 0 164 666 165
rect 0 109 613 164
rect 0 55 666 109
rect 55 54 666 55
rect 55 1 220 54
rect 275 1 385 54
rect 440 1 550 54
rect 605 1 666 54
<< metal2 >>
rect 0 613 118 667
rect 173 613 283 667
rect 338 613 448 667
rect 503 613 613 667
rect 0 604 613 613
rect 0 550 666 604
rect 55 495 666 550
rect 0 494 666 495
rect 0 439 613 494
rect 0 385 666 439
rect 55 330 666 385
rect 0 329 666 330
rect 0 274 613 329
rect 0 220 666 274
rect 55 165 666 220
rect 0 164 666 165
rect 0 109 613 164
rect 0 55 666 109
rect 55 54 666 55
rect 55 1 220 54
rect 275 1 385 54
rect 440 1 550 54
rect 605 1 666 54
<< m123contact >>
rect 118 613 173 667
rect 283 613 338 667
rect 448 613 503 667
rect 613 604 666 667
rect 0 495 55 550
rect 613 439 666 494
rect 0 330 55 385
rect 613 274 666 329
rect 0 165 55 220
rect 613 109 666 164
rect 0 1 55 55
rect 220 1 275 54
rect 385 1 440 54
rect 550 1 605 54
<< metal3 >>
rect 0 613 55 667
rect 173 613 228 667
rect 338 613 393 667
rect 503 613 558 667
rect 0 605 613 613
rect 55 604 613 605
rect 55 549 666 604
rect 55 495 613 549
rect 0 440 613 495
rect 55 439 613 440
rect 55 384 666 439
rect 55 330 613 384
rect 0 275 613 330
rect 55 274 613 275
rect 55 219 666 274
rect 55 165 613 219
rect 0 110 613 165
rect 55 109 613 110
rect 55 54 666 109
rect 165 1 220 54
rect 330 1 385 54
rect 495 1 550 54
<< metal4 >>
rect 118 613 173 667
rect 283 613 338 667
rect 448 613 503 667
rect 613 613 666 667
rect 55 604 666 613
rect 55 550 613 604
rect 0 495 613 550
rect 55 494 613 495
rect 55 439 666 494
rect 55 385 613 439
rect 0 330 613 385
rect 55 329 613 330
rect 55 274 666 329
rect 55 220 613 274
rect 0 165 613 220
rect 55 164 613 165
rect 55 109 666 164
rect 55 55 613 109
rect 0 54 613 55
rect 0 1 55 54
rect 220 1 275 54
rect 385 1 440 54
rect 550 1 605 54
<< m345contact >>
rect 55 613 118 667
rect 228 613 283 667
rect 393 613 448 667
rect 558 613 613 667
rect 0 550 55 605
rect 613 494 666 549
rect 0 385 55 440
rect 613 329 666 384
rect 0 220 55 275
rect 613 164 666 219
rect 0 55 55 110
rect 55 1 165 54
rect 275 1 330 54
rect 440 1 495 54
rect 605 1 666 54
<< metal5 >>
rect 118 613 173 667
rect 283 613 338 667
rect 448 613 503 667
rect 613 613 666 667
rect 55 604 666 613
rect 55 550 613 604
rect 0 495 613 550
rect 55 494 613 495
rect 55 439 666 494
rect 55 385 613 439
rect 0 330 613 385
rect 55 329 613 330
rect 55 274 666 329
rect 55 220 613 274
rect 0 165 613 220
rect 55 164 613 165
rect 55 109 666 164
rect 55 55 613 109
rect 0 54 613 55
rect 0 1 55 54
rect 220 1 275 54
rect 385 1 440 54
rect 550 1 605 54
<< m456contact >>
rect 0 605 55 667
rect 173 613 228 667
rect 338 613 393 667
rect 503 613 558 667
rect 613 549 666 604
rect 0 440 55 495
rect 613 384 666 439
rect 0 275 55 330
rect 613 219 666 274
rect 0 110 55 165
rect 613 54 666 109
rect 165 1 220 54
rect 330 1 385 54
rect 495 1 550 54
<< metal6 >>
rect 55 613 173 667
rect 228 613 338 667
rect 393 613 503 667
rect 558 613 666 667
rect 55 605 666 613
rect 0 604 666 605
rect 0 549 613 604
rect 0 495 666 549
rect 55 440 666 495
rect 0 439 666 440
rect 0 384 613 439
rect 0 330 666 384
rect 55 275 666 330
rect 0 274 666 275
rect 0 219 613 274
rect 0 165 666 219
rect 55 110 666 165
rect 0 109 666 110
rect 0 54 613 109
rect 0 1 165 54
rect 220 1 330 54
rect 385 1 495 54
rect 550 1 666 54
<< glass >>
rect 56 56 612 612
<< end >>
