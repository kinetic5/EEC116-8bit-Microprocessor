magic
tech scmos
timestamp 1575939595
<< error_s >>
rect 97 555 104 558
rect 337 555 344 558
rect 577 555 584 558
rect 817 555 824 558
rect 1057 555 1064 558
rect 1297 555 1304 558
rect 1537 555 1544 558
rect 1777 555 1784 558
rect 104 550 109 551
rect 344 550 349 551
rect 584 550 589 551
rect 824 550 829 551
rect 1064 550 1069 551
rect 1304 550 1309 551
rect 1544 550 1549 551
rect 1784 550 1789 551
rect 101 547 109 550
rect 341 547 349 550
rect 581 547 589 550
rect 821 547 829 550
rect 1061 547 1069 550
rect 1301 547 1309 550
rect 1541 547 1549 550
rect 1781 547 1789 550
rect 233 543 235 546
rect 473 543 475 546
rect 713 543 715 546
rect 953 543 955 546
rect 1193 543 1195 546
rect 1433 543 1435 546
rect 1673 543 1675 546
rect 1913 543 1915 546
rect 53 533 56 543
rect 237 538 239 543
rect 293 533 296 543
rect 477 538 479 543
rect 533 533 536 543
rect 717 538 719 543
rect 773 533 776 543
rect 957 538 959 543
rect 1013 533 1016 543
rect 1197 538 1199 543
rect 1253 533 1256 543
rect 1437 538 1439 543
rect 1493 533 1496 543
rect 1677 538 1679 543
rect 1733 533 1736 543
rect 1917 538 1919 543
rect 1922 542 1923 543
rect 1926 535 1927 542
rect 1922 519 1923 525
rect -133 435 -132 436
rect 275 363 289 364
<< metal1 >>
rect 2141 566 2214 574
rect 2141 506 2185 514
rect 2206 502 2214 566
rect 2141 494 2214 502
rect 2141 434 2185 442
rect 2206 430 2214 494
rect 2141 422 2214 430
rect 2141 362 2185 370
rect 2206 358 2214 422
rect 2141 350 2214 358
rect 2141 290 2185 298
rect 2206 286 2214 350
rect 2141 278 2214 286
rect 2141 218 2185 226
rect 2206 214 2214 278
rect 2141 206 2214 214
rect 2141 146 2185 154
rect 2206 142 2214 206
rect 2141 134 2214 142
rect 2141 74 2185 82
rect 2206 70 2214 134
rect 2141 62 2214 70
rect 2141 2 2185 10
<< m2contact >>
rect 2185 506 2193 514
rect 2185 434 2193 442
rect 2185 362 2193 370
rect 2185 290 2193 298
rect 2185 218 2193 226
rect 2185 146 2193 154
rect 2185 74 2193 82
rect 2185 2 2193 10
<< metal2 >>
rect 37 520 43 524
rect -30 514 43 520
rect -13 441 -7 455
rect 2185 442 2193 506
rect -13 435 73 441
rect 67 427 73 435
rect 227 369 233 383
rect 2185 370 2193 434
rect 227 363 313 369
rect 307 349 313 363
rect 467 297 473 313
rect 2185 298 2193 362
rect 467 291 553 297
rect 547 278 553 291
rect 707 225 713 239
rect 2185 226 2193 290
rect 707 219 793 225
rect 787 206 793 219
rect 947 153 953 168
rect 2185 154 2193 218
rect 947 147 1033 153
rect 1027 133 1033 147
rect 1187 69 1193 95
rect 1147 63 1193 69
rect 2185 82 2193 146
rect 1247 61 1273 67
rect 1247 44 1253 61
rect 2185 10 2193 74
<< m3contact >>
rect -253 543 -247 549
rect 67 471 73 477
rect 307 399 313 405
rect 547 327 553 333
rect 787 255 793 261
rect 1027 183 1033 189
rect 1267 111 1273 117
rect 1507 39 1513 45
<< metal3 >>
rect -243 553 -221 557
rect -95 558 -84 566
rect -287 546 -281 553
rect -243 551 -212 553
rect -247 543 -237 544
rect -297 538 -291 541
rect -253 538 -237 543
rect -228 538 -222 544
rect -218 538 -212 551
rect 12 538 18 552
rect 252 538 258 552
rect 492 538 498 552
rect 732 538 738 552
rect 972 538 978 552
rect 1212 538 1218 552
rect 1452 538 1458 552
rect 1692 538 1698 552
rect 1926 528 1932 542
rect 1937 534 1943 536
rect -87 494 -77 500
rect -83 477 -77 494
rect 225 490 236 494
rect 83 481 99 485
rect 225 486 232 490
rect 33 474 39 481
rect 83 479 108 481
rect 73 471 83 472
rect 23 466 29 469
rect 67 466 83 471
rect 92 464 98 473
rect 102 463 108 479
rect 1925 456 1932 470
rect 1937 462 1943 464
rect 225 429 236 434
rect 157 423 236 429
rect 157 406 163 423
rect 465 419 476 422
rect 323 409 339 413
rect 465 414 477 419
rect 273 402 279 409
rect 323 407 348 409
rect 313 399 329 400
rect 263 394 269 397
rect 307 394 329 399
rect 342 391 348 407
rect 1925 384 1932 398
rect 1937 390 1943 392
rect 387 352 465 357
rect 387 351 476 352
rect 387 333 393 351
rect 563 337 579 341
rect 705 342 716 350
rect 513 330 519 337
rect 563 335 588 337
rect 553 327 569 328
rect 503 322 509 324
rect 547 322 569 327
rect 582 319 588 335
rect 1925 312 1932 326
rect 1937 318 1943 320
rect 705 285 716 290
rect 637 279 716 285
rect 637 261 643 279
rect 803 265 819 269
rect 945 270 956 278
rect 753 258 759 265
rect 803 263 828 265
rect 793 255 809 256
rect 743 250 749 254
rect 787 250 809 255
rect 822 247 828 263
rect 1925 240 1932 254
rect 1937 246 1943 248
rect 945 213 956 218
rect 877 207 956 213
rect 877 190 883 207
rect 1043 193 1059 197
rect 1185 198 1196 206
rect 993 186 999 193
rect 1043 191 1068 193
rect 1033 183 1049 184
rect 983 178 989 181
rect 1027 178 1049 183
rect 1062 173 1068 191
rect 1925 168 1932 182
rect 1937 174 1943 176
rect 1185 141 1196 146
rect 1117 135 1196 141
rect 1117 118 1123 135
rect 1283 121 1299 125
rect 1428 126 1436 134
rect 1233 114 1239 121
rect 1283 119 1308 121
rect 1273 111 1289 112
rect 1223 106 1229 110
rect 1267 106 1289 111
rect 1302 101 1308 119
rect 1925 96 1932 110
rect 1937 102 1943 104
rect 1177 45 1183 62
rect 1357 45 1363 63
rect 1523 49 1539 53
rect 1668 54 1676 62
rect 1473 42 1479 49
rect 1523 47 1548 49
rect 1513 39 1529 40
rect 1463 34 1469 38
rect 1507 34 1529 39
rect 1542 34 1548 47
rect 1897 28 1907 29
rect 1925 28 1932 38
rect 1897 22 1932 28
rect 1937 30 1943 32
<< m4contact >>
rect -95 566 -84 572
rect -182 536 -173 544
rect -122 536 -113 544
rect -74 543 -64 553
rect -55 535 -48 542
rect -13 533 -3 543
rect 101 547 109 554
rect 199 533 207 545
rect 225 538 235 546
rect 341 547 349 554
rect 286 533 296 543
rect 439 533 447 545
rect 465 538 475 546
rect 581 547 589 554
rect 526 533 536 543
rect 679 533 687 545
rect 705 538 715 546
rect 821 547 829 554
rect 766 533 776 543
rect 919 533 927 545
rect 945 538 955 546
rect 1061 547 1069 554
rect 1006 533 1016 543
rect 1159 533 1167 545
rect 1185 538 1195 546
rect 1301 547 1309 554
rect 1246 533 1256 543
rect 1399 533 1407 545
rect 1425 538 1435 546
rect 1541 547 1549 554
rect 1486 533 1496 543
rect 1639 533 1647 545
rect 1665 538 1675 546
rect 1781 547 1789 554
rect 1726 533 1736 543
rect 1879 533 1887 545
rect 1905 538 1915 546
rect 1958 543 1967 550
rect 2077 547 2086 555
rect -96 494 -87 503
rect 225 494 236 500
rect -117 463 -108 472
rect -72 463 -63 472
rect 137 464 147 472
rect 197 464 207 472
rect 406 471 416 481
rect 425 464 435 474
rect 1958 471 1967 478
rect 2077 475 2086 483
rect 225 434 236 440
rect 465 422 476 428
rect 123 391 132 400
rect 168 391 177 400
rect 378 392 387 400
rect 438 392 447 400
rect 646 399 656 409
rect 665 390 675 400
rect 1958 399 1967 406
rect 2077 403 2086 411
rect 465 352 476 358
rect 705 350 716 356
rect 363 319 372 328
rect 410 319 417 328
rect 616 320 627 328
rect 677 320 687 328
rect 887 327 896 336
rect 1958 327 1967 334
rect 2077 331 2086 339
rect 905 318 914 327
rect 705 290 716 296
rect 945 278 956 284
rect 603 246 612 255
rect 648 247 657 256
rect 857 248 867 256
rect 917 248 927 256
rect 1129 255 1136 262
rect 1958 255 1967 262
rect 2077 259 2086 267
rect 1145 245 1155 255
rect 945 218 956 224
rect 1185 206 1196 212
rect 843 174 852 183
rect 888 175 897 184
rect 1097 176 1107 184
rect 1157 176 1167 184
rect 1369 183 1376 190
rect 1385 174 1394 184
rect 1958 183 1967 190
rect 2077 187 2086 195
rect 1185 146 1196 152
rect 1083 103 1092 112
rect 1128 103 1137 112
rect 1336 104 1347 112
rect 1397 104 1407 112
rect 1609 111 1616 118
rect 1625 102 1635 112
rect 1958 111 1967 118
rect 2077 115 2086 123
rect 1177 62 1185 68
rect 1143 31 1152 40
rect 1188 31 1197 40
rect 1323 31 1332 40
rect 1577 32 1587 40
rect 1637 32 1647 40
rect 1849 39 1856 46
rect 1865 30 1874 40
rect 1958 39 1967 46
rect 2077 43 2086 51
<< metal4 >>
rect 225 603 1911 609
rect -195 502 -188 553
rect -182 530 -176 536
rect -150 515 -143 536
rect -120 530 -113 536
rect -95 503 -88 566
rect -83 543 -74 553
rect 102 554 109 578
rect 199 545 207 574
rect -115 472 -108 494
rect -83 3 -76 543
rect -54 530 -48 535
rect 225 546 231 603
rect 342 554 349 578
rect 439 545 447 574
rect 465 546 471 603
rect 582 554 589 578
rect 679 545 687 574
rect 705 546 711 603
rect 822 554 829 578
rect 919 545 927 574
rect 945 546 951 603
rect 1062 554 1069 578
rect 1159 545 1167 574
rect 1185 546 1191 603
rect 1302 554 1309 578
rect 1399 545 1407 574
rect 1425 546 1431 603
rect 1542 554 1549 578
rect 1639 545 1647 574
rect 1665 546 1671 603
rect 1782 554 1789 578
rect 1879 545 1887 574
rect 1905 546 1911 603
rect 2084 578 2085 585
rect 2077 555 2085 578
rect -13 528 -3 533
rect -70 472 -63 504
rect 125 400 132 481
rect 137 451 144 464
rect 170 400 177 464
rect 197 451 204 464
rect 225 440 232 494
rect 289 475 296 533
rect 365 328 372 409
rect 378 380 385 392
rect 399 3 406 481
rect 428 452 435 464
rect 410 328 417 392
rect 440 380 447 392
rect 465 358 472 422
rect 529 403 536 533
rect 634 402 646 409
rect 605 255 612 337
rect 616 308 623 320
rect 634 2 641 402
rect 667 380 675 390
rect 650 256 657 320
rect 680 308 687 320
rect 705 296 712 350
rect 769 331 776 533
rect 876 329 887 336
rect 845 183 852 265
rect 857 236 864 248
rect 876 2 883 329
rect 907 307 914 318
rect 890 184 897 248
rect 920 236 927 248
rect 945 224 952 278
rect 1009 259 1016 533
rect 1115 255 1129 262
rect 1085 112 1092 193
rect 1097 164 1104 176
rect 1115 2 1122 255
rect 1148 236 1155 245
rect 1154 226 1155 236
rect 1130 112 1137 176
rect 1159 164 1167 176
rect 1185 152 1192 206
rect 1249 187 1256 533
rect 1369 151 1376 183
rect 1385 165 1392 174
rect 1145 40 1152 121
rect 1177 68 1184 134
rect 1190 40 1197 104
rect 1336 92 1343 104
rect 1400 92 1407 104
rect 1323 40 1332 49
rect 1412 2 1419 145
rect 1489 115 1496 533
rect 1577 19 1584 32
rect 1609 2 1616 111
rect 1626 92 1633 102
rect 1729 43 1736 533
rect 1639 19 1646 32
rect 1849 3 1856 39
rect 1951 39 1958 550
rect 2077 483 2085 547
rect 2077 411 2085 475
rect 2077 339 2085 403
rect 2077 267 2085 331
rect 2077 195 2085 259
rect 2077 123 2085 187
rect 2077 51 2085 115
rect 1867 20 1874 30
<< m345contact >>
rect -287 553 -278 562
rect -221 553 -212 562
rect -300 529 -291 538
rect -237 536 -228 545
rect 12 552 22 562
rect 46 533 56 543
rect 252 552 262 562
rect 492 552 502 562
rect 732 552 742 562
rect 972 552 982 562
rect 1212 552 1222 562
rect 1452 552 1462 562
rect 1692 552 1702 562
rect 33 481 42 490
rect 99 481 108 490
rect 20 457 29 466
rect 83 464 92 473
rect 273 409 282 418
rect 339 409 348 418
rect 329 394 338 403
rect 260 385 269 394
rect 457 451 467 461
rect 513 337 522 346
rect 579 337 588 346
rect 569 322 578 331
rect 500 313 509 322
rect 697 379 707 389
rect 753 265 762 274
rect 819 265 828 274
rect 809 250 818 259
rect 740 241 749 250
rect 937 307 947 317
rect 993 193 1002 202
rect 1059 193 1068 202
rect 1049 178 1058 187
rect 980 169 989 178
rect 1177 235 1187 245
rect 1417 163 1427 173
rect 1233 121 1242 130
rect 1299 121 1308 130
rect 1289 106 1298 115
rect 1220 97 1229 106
rect 1357 63 1365 69
rect 1368 31 1377 40
rect 1428 134 1436 140
rect 1473 49 1482 58
rect 1539 49 1548 58
rect 1529 34 1538 43
rect 1460 25 1469 34
rect 1657 91 1667 101
rect 1668 62 1676 68
rect 1922 518 1932 528
rect 1937 527 1946 534
rect 1922 446 1932 456
rect 1937 455 1946 462
rect 1922 374 1932 384
rect 1937 383 1946 390
rect 1922 302 1932 312
rect 1937 311 1946 318
rect 1922 230 1932 240
rect 1937 239 1946 246
rect 1922 158 1932 168
rect 1937 167 1946 174
rect 1922 86 1932 96
rect 1937 95 1946 102
rect 1962 527 1971 534
rect 1981 533 1988 545
rect 2128 533 2135 545
rect 1962 455 1971 462
rect 1981 461 1988 473
rect 2128 461 2135 473
rect 1962 383 1971 390
rect 1981 389 1988 401
rect 2128 389 2135 401
rect 1962 311 1971 318
rect 1981 317 1988 329
rect 2128 317 2135 329
rect 1962 239 1971 246
rect 1981 245 1988 257
rect 2128 245 2135 257
rect 1962 167 1971 174
rect 1981 173 1988 185
rect 2128 173 2135 185
rect 1962 95 1971 102
rect 1981 101 1988 113
rect 2128 101 2135 113
rect 1937 23 1946 30
rect 1962 23 1971 30
rect 1981 29 1988 41
rect 2128 29 2135 41
<< m5contact >>
rect 102 578 109 585
rect -197 553 -188 562
rect -152 536 -143 545
rect -182 521 -173 530
rect -122 521 -113 530
rect -150 506 -141 515
rect -195 493 -186 502
rect -117 494 -108 502
rect 342 578 349 585
rect 582 578 589 585
rect 822 578 829 585
rect 1062 578 1069 585
rect 1302 578 1309 585
rect 1542 578 1549 585
rect 1782 578 1789 585
rect 2077 578 2084 585
rect -54 521 -46 530
rect -13 518 -3 528
rect -72 504 -63 513
rect 123 481 132 490
rect 168 464 177 473
rect 137 442 146 451
rect 197 442 206 451
rect 287 466 296 475
rect 363 409 372 418
rect 378 370 388 380
rect 425 442 435 452
rect 410 392 419 401
rect 438 370 448 380
rect 527 394 536 403
rect 603 337 612 346
rect 616 298 626 308
rect -83 -7 -73 3
rect 400 -7 410 3
rect 665 370 675 380
rect 648 320 657 329
rect 677 298 687 308
rect 767 322 776 331
rect 843 265 852 274
rect 857 226 867 236
rect 905 298 914 307
rect 888 248 897 257
rect 917 226 927 236
rect 1007 250 1016 259
rect 1083 193 1092 202
rect 1097 154 1107 164
rect 634 -7 643 2
rect 874 -7 883 2
rect 1144 226 1154 236
rect 1128 176 1137 185
rect 1157 154 1167 164
rect 1247 178 1256 187
rect 1385 155 1396 165
rect 1369 145 1376 151
rect 1412 145 1419 151
rect 1177 134 1185 140
rect 1143 121 1152 130
rect 1188 104 1197 113
rect 1336 82 1346 92
rect 1398 82 1408 92
rect 1323 49 1332 58
rect 1487 106 1496 115
rect 1577 10 1586 19
rect 1623 82 1633 92
rect 1727 34 1736 43
rect 1637 10 1646 19
rect 1866 10 1875 20
rect 1115 -7 1124 2
rect 1412 -7 1421 2
rect 1609 -7 1618 2
rect 1847 -7 1856 3
<< metal5 >>
rect 109 578 342 584
rect 349 578 582 584
rect 589 578 822 584
rect 829 578 1062 584
rect 1069 578 1302 584
rect 1309 578 1542 584
rect 1549 578 1782 584
rect 1789 578 2077 584
rect -320 555 -287 562
rect -278 555 -221 562
rect -212 555 -197 562
rect -188 555 12 562
rect 22 555 252 562
rect 262 555 492 562
rect 502 555 732 562
rect 742 555 972 562
rect 982 555 1212 562
rect 1222 555 1452 562
rect 1462 555 1692 562
rect 1702 555 1913 562
rect -320 538 -237 545
rect -228 538 -152 545
rect -143 543 56 545
rect -143 538 46 543
rect -173 521 -122 527
rect -113 521 -54 527
rect -3 518 1922 525
rect 1946 527 1962 534
rect 1988 533 2128 540
rect -141 506 -72 513
rect -186 494 -117 501
rect -180 483 33 490
rect 42 483 99 490
rect 108 483 123 490
rect 132 483 1920 490
rect -180 466 83 473
rect 92 466 168 473
rect 177 466 287 473
rect 146 442 197 449
rect 206 442 425 449
rect 467 451 1922 453
rect 457 446 1922 451
rect 1946 455 1962 462
rect 1988 461 2128 468
rect 60 411 273 418
rect 282 411 339 418
rect 348 411 363 418
rect 372 411 1913 418
rect 60 394 329 401
rect 338 394 410 401
rect 419 394 527 401
rect 388 370 438 377
rect 448 370 665 377
rect 707 379 1922 381
rect 697 374 1922 379
rect 1946 383 1962 390
rect 1988 389 2128 396
rect 300 339 513 346
rect 522 339 579 346
rect 588 339 603 346
rect 612 339 1913 346
rect 300 322 569 329
rect 578 322 648 329
rect 657 322 767 329
rect 626 298 677 305
rect 947 307 1922 309
rect 687 298 905 305
rect 937 302 1922 307
rect 1946 311 1962 318
rect 1988 317 2128 324
rect 540 267 753 274
rect 762 267 819 274
rect 828 267 843 274
rect 852 267 1913 274
rect 540 250 809 257
rect 818 250 888 257
rect 897 250 1007 257
rect 867 226 917 233
rect 927 226 1144 233
rect 1187 235 1922 237
rect 1177 230 1922 235
rect 1946 239 1962 246
rect 1988 245 2128 252
rect 780 195 993 202
rect 1002 195 1059 202
rect 1068 195 1083 202
rect 1092 195 1913 202
rect 780 178 1049 185
rect 1058 178 1128 185
rect 1137 178 1247 185
rect 1107 154 1157 161
rect 1167 155 1385 162
rect 1427 163 1922 165
rect 1417 158 1922 163
rect 1946 167 1962 174
rect 1988 173 2128 180
rect 1376 145 1412 151
rect 1177 140 1436 141
rect 1185 134 1428 140
rect 1020 123 1143 130
rect 1152 123 1233 130
rect 1242 123 1299 130
rect 1308 123 1913 130
rect 1020 106 1188 113
rect 1197 106 1289 113
rect 1298 106 1487 113
rect 1346 82 1398 89
rect 1408 82 1623 89
rect 1667 91 1922 93
rect 1657 86 1922 91
rect 1946 95 1962 102
rect 1988 101 2128 108
rect 1357 69 1676 70
rect 1365 68 1676 69
rect 1365 63 1668 68
rect 1080 51 1323 58
rect 1332 51 1473 58
rect 1482 51 1539 58
rect 1548 51 1920 58
rect 1260 40 1529 41
rect 1260 34 1368 40
rect 1377 34 1529 40
rect 1538 34 1727 41
rect 1946 23 1962 30
rect 1988 29 2128 36
rect 1586 10 1637 16
rect 1646 10 1866 16
rect -320 -7 -83 0
rect -73 -7 400 0
rect 410 -7 634 0
rect 643 -7 874 0
rect 883 -7 1115 0
rect 1124 -7 1412 0
rect 1421 -7 1609 0
rect 1618 -7 1847 0
rect -320 -18 1920 -11
rect -320 -30 1920 -23
use logic  logic_0
timestamp 1575930433
transform 1 0 -407 0 1 504
box 87 2 327 70
use two_1_mux  two_1_mux_0
timestamp 1575861164
transform 1 0 -125 0 1 565
box 45 -59 125 9
use fadder  fadder_0
timestamp 1575778664
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1575930433
transform 1 0 -87 0 1 432
box 87 2 327 70
use enff  enff_1
timestamp 1575930433
transform 1 0 -269 0 1 362
box -43 -2 148 70
use fadder  fadder_1
timestamp 1575778664
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1575930433
transform 1 0 153 0 1 360
box 87 2 327 70
use enff  enff_2
timestamp 1575930433
transform 1 0 -78 0 1 290
box -43 -2 148 70
use enff  enff_3
timestamp 1575930433
transform 1 0 152 0 1 290
box -43 -2 148 70
use fadder  fadder_2
timestamp 1575778664
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1575930433
transform 1 0 393 0 1 288
box 87 2 327 70
use fadder  fadder_3
timestamp 1575778664
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1575930433
transform 1 0 633 0 1 216
box 87 2 327 70
use fadder  fadder_4
timestamp 1575778664
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1575930433
transform 1 0 873 0 1 144
box 87 2 327 70
use fadder  fadder_5
timestamp 1575778664
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1575930433
transform 1 0 1113 0 1 72
box 87 2 327 70
use fadder  fadder_6
timestamp 1575778664
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1575778664
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1575930433
transform 1 0 1353 0 1 0
box 87 2 327 70
use inv_9_6  inv_9_6_0
array 0 0 30 0 7 72
timestamp 1575933599
transform 1 0 1920 0 1 62
box 0 -60 30 8
use mult  mult_0
timestamp 1575939595
transform 1 0 241 0 1 432
box -241 -432 1689 142
use enff  enff_0
array 0 0 191 0 7 72
timestamp 1575930433
transform 1 0 1993 0 1 2
box -43 -2 148 70
<< labels >>
rlabel m4contact 430 469 430 469 1 4mux_to_2mux_1
rlabel metal4 1884 571 1884 571 1 x7
rlabel metal4 1643 571 1643 571 1 x6
rlabel metal4 1403 570 1403 570 1 x5
rlabel metal4 1163 571 1163 571 1 x4
rlabel metal4 923 570 923 570 1 x3
rlabel metal4 683 570 683 570 1 x2
rlabel metal4 443 570 443 570 1 x1
rlabel metal4 203 570 203 570 1 x0
rlabel metal5 -318 558 -318 558 3 y0
rlabel metal5 -177 486 -177 486 1 y1
rlabel metal5 63 414 63 414 1 y2
rlabel metal5 304 342 304 342 1 y3
rlabel metal5 544 271 544 271 1 y4
rlabel metal5 784 199 784 199 1 y5
rlabel metal5 1025 126 1025 126 1 y6
rlabel metal5 1084 55 1084 55 1 y7
rlabel metal5 -317 -3 -317 -3 3 opcode2
rlabel m5contact 1786 582 1786 582 1 clk
rlabel metal4 1908 605 1908 605 5 x_en
rlabel m4contact -8 535 -8 535 1 nz0
rlabel metal5 1659 88 1659 88 1 nz6
rlabel metal3 1918 25 1918 25 1 nz7
rlabel metal5 459 448 459 448 1 nz1
rlabel m345contact 700 380 700 380 1 nz2
rlabel m345contact 941 308 941 308 1 nz3
rlabel metal5 1181 233 1181 233 1 nz4
rlabel metal5 1420 160 1420 160 1 nz5
rlabel metal5 2123 537 2123 537 1 z0
rlabel metal5 2123 465 2123 465 1 z1
rlabel metal5 2123 392 2123 392 1 z2
rlabel metal5 2123 321 2123 321 1 z3
rlabel metal5 2123 248 2123 248 1 z4
rlabel metal5 2123 176 2123 176 1 z5
rlabel metal5 2123 105 2123 105 1 z6
rlabel metal5 2123 32 2123 32 1 z7
rlabel metal4 1954 546 1954 546 1 c_en
rlabel m2contact 2189 510 2189 510 1 Gnd
rlabel metal1 2210 511 2210 511 7 Vdd
<< end >>
