magic
tech scmos
timestamp 1575998002
<< metal1 >>
rect -3 666 672 668
rect -3 614 58 666
rect 110 614 224 666
rect 279 614 392 666
rect 447 614 560 666
rect 615 614 672 666
rect -3 567 672 614
rect -3 512 -2 567
rect 55 561 672 567
rect 55 512 615 561
rect -3 510 615 512
rect 669 510 672 561
rect -3 405 672 510
rect -3 396 615 405
rect -3 341 -2 396
rect 55 354 615 396
rect 669 354 672 405
rect 55 341 672 354
rect -3 249 672 341
rect -3 225 615 249
rect -3 170 -2 225
rect 55 198 615 225
rect 669 198 672 249
rect 55 170 672 198
rect -3 93 672 170
rect -3 53 615 93
rect -3 52 167 53
rect -3 -3 -2 52
rect 53 -2 167 52
rect 222 -2 335 53
rect 390 -2 503 53
rect 558 42 615 53
rect 669 42 672 93
rect 558 -2 672 42
rect 53 -3 672 -2
rect -3 -4 672 -3
<< metal2 >>
rect -3 666 672 668
rect -3 614 58 666
rect 110 614 224 666
rect 279 614 392 666
rect 447 614 560 666
rect 615 614 672 666
rect -3 567 672 614
rect -3 512 -2 567
rect 55 561 672 567
rect 55 512 615 561
rect -3 510 615 512
rect 669 510 672 561
rect -3 405 672 510
rect -3 396 615 405
rect -3 341 -2 396
rect 55 354 615 396
rect 669 354 672 405
rect 55 341 672 354
rect -3 249 672 341
rect -3 225 615 249
rect -3 170 -2 225
rect 55 198 615 225
rect 669 198 672 249
rect 55 170 672 198
rect -3 93 672 170
rect -3 53 615 93
rect -3 52 167 53
rect -3 -3 -2 52
rect 53 -2 167 52
rect 222 -2 335 53
rect 390 -2 503 53
rect 558 42 615 53
rect 669 42 672 93
rect 558 -2 672 42
rect 53 -3 672 -2
rect -3 -4 672 -3
<< m123contact >>
rect 58 614 110 666
rect 224 614 279 666
rect 392 614 447 666
rect 560 614 615 666
rect -2 512 55 567
rect 615 510 669 561
rect -2 341 55 396
rect 615 354 669 405
rect -2 170 55 225
rect 615 198 669 249
rect -2 -3 53 52
rect 167 -2 222 53
rect 335 -2 390 53
rect 503 -2 558 53
rect 615 42 669 93
<< metal3 >>
rect -3 666 672 668
rect -3 624 58 666
rect -3 569 -2 624
rect 55 614 58 624
rect 110 614 111 666
rect 167 614 224 666
rect 279 614 280 666
rect 335 614 392 666
rect 447 614 448 666
rect 503 614 560 666
rect 615 614 616 666
rect 669 614 672 666
rect 55 569 672 614
rect -3 567 672 569
rect -3 512 -2 567
rect 55 561 672 567
rect 55 512 615 561
rect -3 510 615 512
rect 669 510 672 561
rect -3 509 672 510
rect -3 458 615 509
rect 669 458 672 509
rect -3 453 672 458
rect -3 398 -2 453
rect 55 405 672 453
rect 55 398 615 405
rect -3 396 615 398
rect -3 341 -2 396
rect 55 354 615 396
rect 669 354 672 405
rect 55 353 672 354
rect 55 341 615 353
rect -3 302 615 341
rect 669 302 672 353
rect -3 282 672 302
rect -3 227 -2 282
rect 55 249 672 282
rect 55 227 615 249
rect -3 225 615 227
rect -3 170 -2 225
rect 55 198 615 225
rect 669 198 672 249
rect 55 197 672 198
rect 55 170 615 197
rect -3 147 615 170
rect 669 147 672 197
rect -3 111 672 147
rect -3 54 -2 111
rect 55 93 672 111
rect 55 54 615 93
rect -3 53 615 54
rect -3 52 111 53
rect -3 -3 -2 52
rect 53 -2 111 52
rect 166 -2 167 53
rect 222 -2 279 53
rect 334 -2 335 53
rect 390 -2 447 53
rect 502 -2 503 53
rect 558 42 615 53
rect 669 42 672 93
rect 558 40 672 42
rect 558 -2 615 40
rect 669 -2 672 40
rect 53 -3 672 -2
rect -3 -4 672 -3
<< metal4 >>
rect -3 667 672 668
rect -3 626 -2 667
rect 55 666 672 667
rect 55 626 111 666
rect -3 624 111 626
rect -3 569 -2 624
rect 55 614 111 624
rect 167 614 168 666
rect 223 614 280 666
rect 335 614 336 666
rect 391 614 448 666
rect 503 614 504 666
rect 559 614 616 666
rect 669 614 672 666
rect 55 613 672 614
rect 55 569 615 613
rect -3 562 615 569
rect 669 562 672 613
rect -3 510 672 562
rect -3 455 -2 510
rect 55 509 672 510
rect 55 458 615 509
rect 669 458 672 509
rect 55 457 672 458
rect 55 455 615 457
rect -3 453 615 455
rect -3 398 -2 453
rect 55 406 615 453
rect 669 406 672 457
rect 55 398 672 406
rect -3 353 672 398
rect -3 339 615 353
rect -3 284 -2 339
rect 55 302 615 339
rect 669 302 672 353
rect 55 301 672 302
rect 55 284 615 301
rect -3 282 615 284
rect -3 227 -2 282
rect 55 250 615 282
rect 669 250 672 301
rect 55 227 672 250
rect -3 197 672 227
rect -3 168 615 197
rect -3 113 -2 168
rect 55 147 615 168
rect 669 147 672 197
rect 55 145 672 147
rect 55 113 615 145
rect -3 111 615 113
rect -3 54 -2 111
rect 55 94 615 111
rect 669 94 672 145
rect 55 54 672 94
rect -3 53 672 54
rect -3 -2 55 53
rect 110 -2 111 53
rect 166 -2 223 53
rect 278 -2 279 53
rect 334 -2 391 53
rect 446 -2 447 53
rect 502 -2 559 53
rect 614 40 672 53
rect 614 -2 615 40
rect 669 -2 672 40
rect -3 -4 672 -2
<< m345contact >>
rect -2 569 55 624
rect 111 614 167 666
rect 280 614 335 666
rect 448 614 503 666
rect 616 614 669 666
rect 615 458 669 509
rect -2 398 55 453
rect 615 302 669 353
rect -2 227 55 282
rect 615 147 669 197
rect -2 54 55 111
rect 111 -2 166 53
rect 279 -2 334 53
rect 447 -2 502 53
rect 615 -2 669 40
<< metal5 >>
rect -3 667 672 668
rect -3 626 -2 667
rect 55 666 672 667
rect 55 626 111 666
rect -3 624 111 626
rect -3 569 -2 624
rect 55 614 111 624
rect 167 614 168 666
rect 223 614 280 666
rect 335 614 336 666
rect 391 614 448 666
rect 503 614 504 666
rect 559 614 616 666
rect 669 614 672 666
rect 55 613 672 614
rect 55 569 615 613
rect -3 562 615 569
rect 669 562 672 613
rect -3 510 672 562
rect -3 455 -2 510
rect 55 509 672 510
rect 55 458 615 509
rect 669 458 672 509
rect 55 457 672 458
rect 55 455 615 457
rect -3 453 615 455
rect -3 398 -2 453
rect 55 406 615 453
rect 669 406 672 457
rect 55 398 672 406
rect -3 353 672 398
rect -3 339 615 353
rect -3 284 -2 339
rect 55 302 615 339
rect 669 302 672 353
rect 55 301 672 302
rect 55 284 615 301
rect -3 282 615 284
rect -3 227 -2 282
rect 55 250 615 282
rect 669 250 672 301
rect 55 227 672 250
rect -3 197 672 227
rect -3 168 615 197
rect -3 113 -2 168
rect 55 147 615 168
rect 669 147 672 197
rect 55 145 672 147
rect 55 113 615 145
rect -3 111 615 113
rect -3 54 -2 111
rect 55 94 615 111
rect 669 94 672 145
rect 55 54 672 94
rect -3 53 672 54
rect -3 -2 55 53
rect 110 -2 111 53
rect 166 -2 223 53
rect 278 -2 279 53
rect 334 -2 391 53
rect 446 -2 447 53
rect 502 -2 559 53
rect 614 40 672 53
rect 614 -2 615 40
rect 669 -2 672 40
rect -3 -4 672 -2
<< m456contact >>
rect -2 626 55 667
rect 168 614 223 666
rect 336 614 391 666
rect 504 614 559 666
rect 615 562 669 613
rect -2 455 55 510
rect 615 406 669 457
rect -2 284 55 339
rect 615 250 669 301
rect -2 113 55 168
rect 615 94 669 145
rect 55 -2 110 53
rect 223 -2 278 53
rect 391 -2 446 53
rect 559 -2 614 53
<< metal6 >>
rect -3 667 672 668
rect -3 626 -2 667
rect 55 666 672 667
rect 55 626 168 666
rect -3 614 168 626
rect 223 614 336 666
rect 391 614 504 666
rect 559 614 672 666
rect -3 613 672 614
rect -3 562 615 613
rect 669 562 672 613
rect -3 510 672 562
rect -3 455 -2 510
rect 55 457 672 510
rect 55 455 615 457
rect -3 406 615 455
rect 669 406 672 457
rect -3 339 672 406
rect -3 284 -2 339
rect 55 301 672 339
rect 55 284 615 301
rect -3 250 615 284
rect 669 250 672 301
rect -3 168 672 250
rect -3 113 -2 168
rect 55 145 672 168
rect 55 113 615 145
rect -3 94 615 113
rect 669 94 672 145
rect -3 53 672 94
rect -3 -2 55 53
rect 110 -2 223 53
rect 278 -2 391 53
rect 446 -2 559 53
rect 614 -2 672 53
rect -3 -4 672 -2
<< glass >>
rect 56 56 612 612
<< end >>
