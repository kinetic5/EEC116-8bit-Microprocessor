magic
tech scmos
timestamp 1575960871
<< metal1 >>
rect 2138 566 2214 574
rect 2137 506 2185 514
rect 2206 502 2214 566
rect 2140 494 2214 502
rect 2136 434 2185 442
rect 2206 430 2214 494
rect 2138 422 2214 430
rect 2138 362 2185 370
rect 2206 358 2214 422
rect 2138 350 2214 358
rect 2136 290 2185 298
rect 2206 286 2214 350
rect 2135 278 2214 286
rect 2138 218 2185 226
rect 2206 214 2214 278
rect 2139 206 2214 214
rect 2139 146 2185 154
rect 2206 142 2214 206
rect 2139 134 2214 142
rect 2137 74 2185 82
rect 2206 70 2214 134
rect 2137 62 2214 70
rect 2138 2 2185 10
<< m2contact >>
rect 2185 506 2193 514
rect 2185 434 2193 442
rect 2185 362 2193 370
rect 2185 290 2193 298
rect 2185 218 2193 226
rect 2185 146 2193 154
rect 2185 74 2193 82
rect 2185 2 2193 10
<< metal2 >>
rect 37 520 43 524
rect -30 514 43 520
rect -213 505 -208 506
rect -13 441 -7 455
rect 2185 442 2193 506
rect -13 435 73 441
rect 67 427 73 435
rect 107 431 144 436
rect 139 429 144 431
rect 139 424 148 429
rect 227 369 233 383
rect 2185 370 2193 434
rect 227 363 313 369
rect 307 349 313 363
rect 347 359 383 365
rect 377 358 383 359
rect 467 297 473 313
rect 2185 298 2193 362
rect 467 291 553 297
rect 547 278 553 291
rect 587 288 624 292
rect 620 279 624 288
rect 707 225 713 239
rect 2185 226 2193 290
rect 707 219 793 225
rect 787 206 793 219
rect 827 217 862 221
rect 859 207 863 217
rect 947 153 953 168
rect 2185 154 2193 218
rect 947 147 1033 153
rect 1027 133 1033 147
rect 1067 143 1105 148
rect 1100 135 1105 143
rect 1187 69 1193 95
rect 2185 82 2193 146
rect 1279 75 1312 76
rect 1279 74 1307 75
rect 1238 72 1312 74
rect 1147 63 1193 69
rect 1236 71 1312 72
rect 1236 69 1242 71
rect 1307 70 1312 71
rect 1247 61 1273 67
rect 1247 44 1253 61
rect 2185 10 2193 74
<< m3contact >>
rect -253 543 -247 549
rect -213 500 -208 505
rect 67 471 73 477
rect 148 424 154 430
rect 307 399 313 405
rect 377 352 383 358
rect 547 327 553 333
rect 624 279 630 285
rect 787 255 793 261
rect 863 207 869 213
rect 1027 183 1033 189
rect 1105 135 1111 141
rect 1267 111 1273 117
rect 1236 63 1242 69
rect 1507 39 1513 45
<< metal3 >>
rect -243 553 -222 557
rect -95 558 -84 566
rect -287 546 -281 553
rect -243 551 -212 553
rect -247 543 -237 544
rect -297 538 -291 541
rect -253 538 -237 543
rect -228 538 -222 544
rect -218 538 -212 551
rect 12 538 18 552
rect 252 538 258 552
rect 492 538 498 552
rect 732 538 738 552
rect 972 538 978 552
rect 1212 538 1218 552
rect 1452 538 1458 552
rect 1692 538 1698 552
rect 1927 528 1933 542
rect 1943 536 1945 542
rect 1937 534 1947 536
rect 1970 527 1975 531
rect 225 490 236 494
rect 83 481 98 485
rect 225 486 232 490
rect 33 474 39 481
rect 83 479 108 481
rect 73 471 83 472
rect 23 466 29 469
rect 67 466 83 471
rect 92 464 98 473
rect 102 463 108 479
rect 457 457 467 461
rect 1925 456 1932 470
rect 1937 462 1943 464
rect 1970 455 1975 460
rect 154 424 163 430
rect 157 406 163 424
rect 465 419 476 422
rect 323 409 338 413
rect 465 414 477 419
rect 273 402 279 409
rect 323 407 348 409
rect -53 389 -34 401
rect 313 399 329 400
rect 263 394 269 397
rect 307 394 329 399
rect 342 391 348 407
rect 1925 384 1932 398
rect 1937 390 1943 392
rect 1970 383 1975 387
rect 383 352 393 358
rect 387 333 393 352
rect 563 337 578 341
rect 705 342 716 350
rect 513 330 519 337
rect 563 335 588 337
rect -123 317 -104 329
rect 187 317 206 329
rect 553 327 569 328
rect 503 322 509 324
rect 547 322 569 327
rect 582 319 588 335
rect 1925 312 1932 326
rect 1937 318 1943 320
rect 1970 311 1975 315
rect 690 285 698 290
rect 630 279 643 285
rect 637 261 643 279
rect 803 265 818 269
rect 945 270 956 278
rect 753 258 759 265
rect 803 263 828 265
rect -320 247 -313 255
rect -177 240 -174 258
rect -126 246 -95 256
rect 117 245 136 257
rect 427 245 446 257
rect 793 255 809 256
rect 743 250 749 254
rect 787 250 809 255
rect 822 247 828 263
rect 1925 240 1932 254
rect 1937 246 1943 248
rect 1970 239 1975 243
rect 869 207 883 213
rect 877 190 883 207
rect 1043 193 1058 197
rect 1185 198 1196 206
rect 993 186 999 193
rect 1043 191 1068 193
rect -107 168 -104 186
rect 133 168 136 186
rect 373 168 376 186
rect 667 173 686 185
rect 1033 183 1049 184
rect 983 178 989 181
rect 1027 178 1049 183
rect 1062 173 1068 191
rect 1925 168 1932 182
rect 1937 174 1943 176
rect 1970 167 1975 171
rect 1111 135 1123 141
rect 1117 118 1123 135
rect 1283 121 1298 125
rect 1428 126 1436 134
rect 1233 114 1239 121
rect 1283 119 1308 121
rect 907 101 926 113
rect 1273 111 1289 112
rect 1223 106 1229 110
rect 1267 106 1289 111
rect 1302 101 1308 119
rect 1925 96 1932 110
rect 1937 102 1943 104
rect 1970 95 1975 99
rect 1177 63 1236 69
rect 1242 63 1244 69
rect 1177 45 1183 63
rect 1357 45 1363 63
rect 1523 49 1538 53
rect 1668 54 1676 62
rect 1473 42 1479 49
rect 1523 47 1548 49
rect 967 29 986 41
rect 1513 39 1529 40
rect 1463 34 1469 38
rect 1507 34 1529 39
rect 1542 34 1548 47
rect 1897 28 1907 29
rect 1925 28 1932 38
rect 1897 22 1932 28
rect 1937 30 1943 32
rect 1970 23 1975 27
<< m4contact >>
rect -178 568 -170 574
rect -150 568 -142 574
rect -106 568 -99 574
rect -95 566 -84 572
rect -208 545 -202 553
rect -182 536 -173 544
rect -122 536 -113 544
rect -74 543 -64 553
rect -55 535 -48 542
rect -13 533 -3 543
rect 109 546 119 554
rect 139 547 147 554
rect 235 543 243 555
rect 349 546 359 554
rect 379 547 387 554
rect 475 543 483 555
rect 283 533 293 543
rect 589 546 599 554
rect 619 547 627 554
rect 715 543 723 555
rect 523 533 533 543
rect 829 546 839 554
rect 859 547 867 554
rect 955 543 963 555
rect 763 533 773 543
rect 1069 546 1079 554
rect 1099 547 1107 554
rect 1195 543 1203 555
rect 1003 533 1013 543
rect 1309 546 1319 554
rect 1339 547 1347 554
rect 1435 543 1443 555
rect 1243 533 1253 543
rect 1549 546 1559 554
rect 1579 547 1587 554
rect 1675 543 1683 555
rect 1483 533 1493 543
rect 1789 546 1799 554
rect 1819 547 1827 554
rect 1915 543 1923 555
rect 1957 543 1966 550
rect 2076 547 2085 555
rect 1723 533 1733 543
rect -178 506 -170 512
rect -110 506 -102 512
rect 142 496 150 502
rect 179 496 190 502
rect 210 496 221 502
rect -117 463 -108 472
rect -72 463 -63 472
rect 113 475 118 483
rect 137 464 147 472
rect 197 464 207 472
rect 406 471 416 481
rect 425 464 435 474
rect 1957 471 1966 478
rect 2076 475 2085 483
rect 138 434 150 440
rect 210 434 222 440
rect 192 426 198 434
rect 384 424 390 430
rect 422 424 430 430
rect 450 424 458 430
rect 45 390 55 400
rect 123 391 132 400
rect 168 391 177 400
rect 352 403 358 409
rect 378 392 387 400
rect 438 392 447 400
rect 646 399 656 409
rect 665 390 675 400
rect 1957 399 1966 406
rect 2076 403 2085 411
rect 422 360 429 366
rect 622 352 630 357
rect 650 352 658 358
rect 690 352 698 357
rect -25 318 -15 328
rect 285 318 295 328
rect 363 319 372 328
rect 410 319 417 328
rect 592 331 598 337
rect 616 320 627 328
rect 677 320 687 328
rect 887 327 896 336
rect 1957 327 1966 334
rect 2076 331 2085 339
rect 905 318 914 327
rect 662 285 670 291
rect 862 280 870 286
rect 902 280 910 286
rect 930 280 938 286
rect -136 246 -126 256
rect 215 246 225 256
rect 525 246 535 256
rect 603 246 612 255
rect 648 247 657 256
rect 832 258 838 264
rect 857 248 867 256
rect 920 248 927 256
rect 1129 255 1136 262
rect 1957 255 1966 262
rect 2076 259 2085 267
rect 1145 245 1155 255
rect 862 217 870 222
rect 901 218 907 224
rect 1102 208 1110 214
rect 1141 208 1150 214
rect 1170 208 1179 214
rect -250 171 -243 183
rect -10 171 -3 183
rect 230 171 237 183
rect 765 174 775 184
rect 843 174 852 183
rect 888 175 897 184
rect 1072 186 1078 193
rect 1097 176 1107 184
rect 1157 176 1167 184
rect 1369 183 1376 190
rect 1385 174 1394 184
rect 1957 183 1966 190
rect 2076 187 2085 195
rect 1102 145 1110 150
rect 1142 146 1150 152
rect 1171 146 1179 152
rect 1342 136 1348 142
rect 1378 136 1390 142
rect 1402 126 1408 136
rect 1005 102 1015 112
rect 1083 103 1092 112
rect 1128 103 1137 112
rect 1312 114 1318 121
rect 1336 104 1347 112
rect 1397 104 1407 112
rect 1609 111 1616 118
rect 1625 102 1635 112
rect 1957 111 1966 118
rect 2076 115 2085 123
rect 1347 66 1353 74
rect 1392 66 1398 74
rect 1402 66 1408 74
rect 1582 64 1590 70
rect 1622 64 1630 70
rect 1650 64 1658 70
rect 1065 30 1075 40
rect 1143 31 1152 40
rect 1188 31 1197 40
rect 1323 31 1332 40
rect 1577 32 1587 40
rect 1637 32 1647 40
rect 1849 39 1856 46
rect 1865 30 1874 40
rect 1957 39 1966 46
rect 2076 43 2085 51
rect 1650 2 1658 8
rect 1590 -4 1598 2
rect 1630 -4 1638 2
<< metal4 >>
rect -208 553 -202 578
rect -206 462 -199 496
rect -195 502 -188 553
rect -182 530 -176 536
rect -150 515 -143 536
rect -136 256 -129 566
rect -117 564 -110 584
rect -90 572 -84 578
rect -117 557 -102 564
rect -120 530 -113 536
rect -109 512 -102 557
rect -94 546 -74 553
rect -110 472 -103 494
rect -108 463 -103 472
rect -94 214 -87 546
rect -76 543 -74 546
rect -54 530 -48 535
rect -13 528 -3 533
rect -70 472 -63 504
rect -25 328 -18 481
rect 58 400 65 552
rect 109 554 115 567
rect 140 554 147 578
rect 235 555 243 584
rect 349 554 355 567
rect 380 554 387 578
rect 475 555 483 584
rect 589 554 596 567
rect 620 554 627 578
rect 715 555 721 596
rect 829 554 835 567
rect 860 554 867 578
rect 955 555 963 589
rect 1069 554 1075 567
rect 1100 554 1107 578
rect 1195 555 1203 584
rect 1309 554 1315 567
rect 1340 554 1347 578
rect 1435 555 1443 584
rect 1549 554 1555 567
rect 1580 554 1587 578
rect 1675 555 1683 584
rect 1793 554 1799 567
rect 1820 554 1827 578
rect 1915 555 1923 584
rect 2084 578 2085 585
rect 2077 555 2085 578
rect 1951 543 1957 550
rect 142 502 149 505
rect 113 483 117 495
rect 125 400 132 481
rect 137 453 144 464
rect 157 440 164 506
rect 210 502 217 506
rect 150 433 164 440
rect 55 390 65 400
rect -250 -74 -243 171
rect -10 -74 -3 171
rect 157 2 164 433
rect 170 400 177 466
rect 181 2 188 496
rect 286 475 293 533
rect 197 449 204 464
rect 192 3 198 426
rect 210 429 218 434
rect 384 430 390 460
rect 352 409 358 424
rect 218 256 225 337
rect 288 328 295 409
rect 365 328 372 409
rect 378 382 385 392
rect 230 -74 237 171
rect 383 1 390 362
rect 399 3 406 481
rect 428 452 435 464
rect 452 434 458 442
rect 450 430 458 434
rect 410 328 417 392
rect 424 376 430 424
rect 440 387 447 392
rect 440 380 450 387
rect 424 370 438 376
rect 422 2 429 360
rect 433 364 438 370
rect 433 2 439 364
rect 480 362 486 460
rect 526 403 533 533
rect 634 402 646 409
rect 451 0 458 356
rect 592 337 597 352
rect 620 357 625 358
rect 620 352 622 357
rect 528 256 535 264
rect 605 255 612 337
rect 616 308 623 320
rect 623 2 630 289
rect 634 2 641 402
rect 650 358 658 381
rect 667 380 675 390
rect 698 352 701 357
rect 650 256 657 320
rect 680 308 687 320
rect 694 294 701 352
rect 766 331 773 533
rect 876 329 887 336
rect 662 2 669 285
rect 833 264 837 278
rect 768 184 775 193
rect 845 183 852 265
rect 857 236 864 248
rect 876 2 883 329
rect 907 307 914 318
rect 910 280 916 286
rect 890 184 897 248
rect 901 2 907 218
rect 911 2 916 280
rect 920 236 927 248
rect 931 231 936 280
rect 931 226 947 231
rect 942 212 947 226
rect 942 2 947 207
rect 960 222 966 288
rect 1006 259 1013 533
rect 1115 255 1129 262
rect 960 2 966 216
rect 1072 193 1077 206
rect 1008 112 1015 120
rect 1085 112 1092 193
rect 1097 164 1104 176
rect 1068 40 1075 49
rect 1103 0 1109 145
rect 1115 2 1122 255
rect 1148 236 1155 245
rect 1154 226 1155 236
rect 1246 187 1253 533
rect 1130 112 1137 176
rect 1159 164 1167 176
rect 1369 151 1376 183
rect 1385 165 1392 174
rect 1142 140 1148 146
rect 1142 134 1162 140
rect 1145 40 1152 121
rect 1156 1 1162 134
rect 1170 1 1176 146
rect 1374 146 1376 151
rect 1342 142 1348 143
rect 1312 121 1317 134
rect 1190 40 1197 104
rect 1336 92 1343 104
rect 1347 74 1353 94
rect 1323 40 1332 49
rect 1335 -11 1341 4
rect 1347 -34 1353 66
rect 1378 50 1384 136
rect 1402 124 1408 126
rect 1388 118 1408 124
rect 1388 102 1393 118
rect 1400 92 1407 104
rect 1378 44 1387 50
rect 1381 -45 1387 44
rect 1392 -23 1398 66
rect 1402 -12 1408 66
rect 1412 2 1419 145
rect 1486 115 1493 533
rect 1567 64 1582 70
rect 1567 -11 1573 64
rect 1577 16 1584 32
rect 1609 2 1616 111
rect 1626 92 1633 102
rect 1590 -33 1597 -4
rect 1620 64 1622 70
rect 1658 64 1664 70
rect 1620 -22 1626 64
rect 1639 16 1646 32
rect 1657 19 1664 64
rect 1726 43 1733 533
rect 1951 478 1958 543
rect 2077 483 2085 547
rect 1951 471 1957 478
rect 1951 406 1958 471
rect 2077 411 2085 475
rect 1951 399 1957 406
rect 1951 334 1958 399
rect 2077 339 2085 403
rect 1951 327 1957 334
rect 1951 262 1958 327
rect 2077 267 2085 331
rect 1951 255 1957 262
rect 1951 190 1958 255
rect 2077 195 2085 259
rect 1951 183 1957 190
rect 1951 118 1958 183
rect 2077 123 2085 187
rect 1951 111 1957 118
rect 1951 46 1958 111
rect 2077 51 2085 115
rect 1657 12 1669 19
rect 1630 -44 1637 -4
rect 1650 -11 1657 2
rect 1662 -33 1669 12
rect 1849 3 1856 39
rect 1951 39 1957 46
rect 1867 20 1874 30
<< m345contact >>
rect -287 553 -278 562
rect -222 553 -213 562
rect -300 529 -291 538
rect -237 536 -228 545
rect -208 496 -199 505
rect 12 552 22 562
rect 43 533 53 543
rect 33 481 42 490
rect -83 453 -76 461
rect 20 457 29 466
rect 252 552 262 562
rect 492 552 502 562
rect 732 552 742 562
rect 972 552 982 562
rect 1212 552 1222 562
rect 1452 552 1462 562
rect 1692 552 1702 562
rect 98 481 107 490
rect 83 464 92 473
rect 225 494 236 500
rect 273 409 282 418
rect 338 409 347 418
rect 260 385 269 394
rect 329 394 338 403
rect 382 362 390 368
rect 457 447 467 457
rect 465 422 476 428
rect 450 356 458 362
rect 513 337 522 346
rect 578 337 587 346
rect 569 322 578 331
rect 500 313 509 322
rect 622 289 630 294
rect 697 379 707 389
rect 705 350 716 356
rect 690 279 698 285
rect 753 265 762 274
rect 818 265 827 274
rect 809 250 818 259
rect 740 241 749 250
rect 937 307 947 317
rect 945 278 956 284
rect 930 216 938 222
rect 993 193 1002 202
rect 1058 193 1067 202
rect 1049 178 1058 187
rect 980 169 989 178
rect 1177 235 1187 245
rect 1185 206 1196 212
rect 1417 163 1427 173
rect 1233 121 1242 130
rect 1298 121 1307 130
rect 1289 106 1298 115
rect 1220 97 1229 106
rect 1357 63 1365 69
rect 1368 31 1377 40
rect 1428 134 1436 140
rect 1473 49 1482 58
rect 1538 49 1547 58
rect 1529 34 1538 43
rect 1460 25 1469 34
rect 1657 91 1667 101
rect 1668 62 1676 68
rect 1927 518 1934 528
rect 1938 527 1947 534
rect 1962 527 1970 534
rect 1980 533 1987 545
rect 2128 533 2135 545
rect 1922 446 1932 456
rect 1937 455 1946 462
rect 1962 455 1970 462
rect 1980 461 1987 473
rect 2128 461 2135 473
rect 1922 374 1932 384
rect 1937 383 1946 390
rect 1962 383 1970 390
rect 1980 389 1987 401
rect 2128 389 2135 401
rect 1922 302 1932 312
rect 1937 311 1946 318
rect 1962 311 1970 318
rect 1980 317 1987 329
rect 2128 317 2135 329
rect 1922 230 1932 240
rect 1937 239 1946 246
rect 1962 239 1970 246
rect 1980 245 1987 257
rect 2128 245 2135 257
rect 1922 158 1932 168
rect 1937 167 1946 174
rect 1962 167 1970 174
rect 1980 173 1987 185
rect 2128 173 2135 185
rect 1922 86 1932 96
rect 1937 95 1946 102
rect 1962 95 1970 102
rect 1980 101 1987 113
rect 2128 101 2135 113
rect 1937 23 1946 30
rect 1962 23 1970 30
rect 1980 29 1987 41
rect 2128 29 2135 41
<< m5contact >>
rect -208 578 -202 584
rect -136 566 -121 574
rect -197 553 -188 562
rect -152 536 -143 545
rect -182 521 -173 530
rect -150 506 -141 515
rect -195 493 -186 502
rect -206 453 -197 462
rect -90 578 -84 584
rect 140 578 147 585
rect 109 567 116 574
rect -122 521 -113 530
rect -112 494 -103 502
rect 55 552 65 562
rect -54 521 -46 530
rect -13 518 -3 528
rect -72 504 -63 513
rect -27 481 -18 490
rect 380 578 387 585
rect 349 567 356 574
rect 620 578 627 584
rect 589 567 596 574
rect 860 578 867 585
rect 829 567 836 574
rect 1100 578 1107 585
rect 1069 567 1076 574
rect 1340 578 1347 585
rect 1309 567 1316 574
rect 1580 578 1587 585
rect 1549 567 1556 574
rect 1820 578 1827 585
rect 1793 567 1800 574
rect 2077 578 2084 585
rect 157 506 164 513
rect 113 495 119 501
rect 123 481 132 490
rect 137 444 146 453
rect 210 506 217 513
rect 168 466 177 473
rect -83 -7 -73 3
rect 284 466 293 475
rect 384 460 390 466
rect 197 442 206 449
rect 210 422 218 429
rect 352 424 358 430
rect 286 409 295 418
rect 363 409 372 418
rect 216 337 225 346
rect 378 372 388 382
rect 480 460 486 466
rect 425 442 435 452
rect 410 392 419 401
rect 442 370 450 380
rect 400 -7 410 3
rect 524 394 533 403
rect 478 356 486 362
rect 592 352 599 358
rect 603 337 612 346
rect 528 264 538 274
rect 616 298 626 308
rect 665 370 675 380
rect 648 320 657 329
rect 677 298 687 308
rect 764 322 773 331
rect 694 289 701 294
rect 862 286 871 292
rect 833 278 840 284
rect 843 265 852 274
rect 768 193 777 202
rect 857 226 867 236
rect 862 212 870 217
rect 905 298 914 307
rect 960 288 966 294
rect 888 248 897 257
rect 920 226 927 236
rect 942 207 947 212
rect 1004 250 1013 259
rect 960 216 966 222
rect 1072 206 1080 212
rect 1083 193 1092 202
rect 1008 120 1018 130
rect 1097 154 1107 164
rect 1068 49 1077 58
rect 634 -7 643 2
rect 874 -7 883 2
rect 1144 226 1154 236
rect 1128 176 1137 185
rect 1244 178 1253 187
rect 1157 154 1167 164
rect 1385 155 1396 165
rect 1143 121 1152 130
rect 1115 -7 1124 2
rect 1368 145 1374 151
rect 1412 145 1419 151
rect 1312 134 1319 141
rect 1188 104 1197 113
rect 1336 82 1343 92
rect 1347 94 1353 100
rect 1323 49 1332 58
rect 1335 -18 1341 -11
rect 1388 95 1393 102
rect 1398 82 1408 92
rect 1347 -40 1353 -34
rect 1484 106 1493 115
rect 1412 -7 1421 2
rect 1402 -18 1408 -12
rect 1577 10 1586 16
rect 1623 82 1633 92
rect 1567 -18 1574 -11
rect 1392 -29 1398 -23
rect 1607 -7 1616 2
rect 1637 10 1646 16
rect 1724 34 1733 43
rect 1618 -29 1626 -22
rect 1590 -40 1598 -33
rect 1381 -51 1387 -45
rect 1650 -18 1658 -11
rect 1866 10 1875 20
rect 1847 -7 1856 3
rect 1662 -40 1670 -33
rect 1630 -51 1638 -44
<< metal5 >>
rect -202 578 -90 584
rect 109 578 140 584
rect 147 578 380 584
rect 387 578 620 584
rect 627 578 860 584
rect 867 578 1100 584
rect 1107 578 1340 584
rect 1347 578 1580 584
rect 1587 578 1820 584
rect 1827 578 2077 584
rect -121 567 109 574
rect 116 567 349 574
rect 356 567 589 574
rect 596 567 829 574
rect 836 567 1069 574
rect 1076 567 1309 574
rect 1316 567 1549 574
rect 1556 567 1793 574
rect -320 555 -287 562
rect -278 555 -222 562
rect -213 555 -197 562
rect -188 555 12 562
rect 22 555 55 562
rect 65 555 252 562
rect 262 555 492 562
rect 502 555 732 562
rect 742 555 972 562
rect 982 555 1212 562
rect 1222 555 1452 562
rect 1462 555 1692 562
rect 1702 555 1913 562
rect -320 538 -237 545
rect -228 538 -152 545
rect -143 543 53 545
rect -143 538 43 543
rect -173 521 -122 527
rect -113 521 -54 527
rect -3 518 1927 525
rect 1947 527 1962 534
rect 1987 533 2128 540
rect -141 506 -72 513
rect 164 507 210 513
rect -186 494 -112 501
rect 119 495 225 500
rect -180 483 -27 490
rect -18 483 33 490
rect 42 483 98 490
rect 107 483 123 490
rect 132 483 1920 490
rect -180 466 83 473
rect -197 453 -83 460
rect 92 466 168 473
rect 177 466 284 473
rect 447 466 471 467
rect 390 461 480 466
rect 390 460 453 461
rect 471 460 480 461
rect 146 444 197 449
rect 137 442 197 444
rect 206 442 425 449
rect 467 447 1922 453
rect 457 446 1922 447
rect 1946 455 1962 462
rect 1987 461 2128 468
rect 149 422 210 429
rect 358 428 476 430
rect 358 424 465 428
rect 60 411 273 418
rect 282 411 286 418
rect 295 411 338 418
rect 348 411 363 418
rect 372 411 1913 418
rect 60 394 329 401
rect 338 394 410 401
rect 419 394 524 401
rect 388 372 442 377
rect 394 370 442 372
rect 450 370 665 377
rect 707 379 1922 381
rect 697 374 1922 379
rect 1946 383 1962 390
rect 1987 389 2128 396
rect 592 362 716 366
rect 458 356 478 362
rect 592 361 601 362
rect 624 361 716 362
rect 592 358 599 361
rect 705 356 716 361
rect 225 339 513 346
rect 522 339 578 346
rect 587 339 603 346
rect 612 339 1913 346
rect 300 322 569 329
rect 578 322 648 329
rect 657 322 764 329
rect 626 298 677 305
rect 947 307 1922 309
rect 687 298 905 305
rect 937 302 1922 307
rect 1946 311 1962 318
rect 1987 317 2128 324
rect 630 289 694 294
rect 862 292 960 294
rect 871 288 960 292
rect 618 279 690 284
rect 618 278 698 279
rect 840 278 945 282
rect 538 267 753 274
rect 762 267 818 274
rect 828 267 843 274
rect 852 267 1913 274
rect 540 250 809 257
rect 818 250 888 257
rect 897 250 1004 257
rect 867 226 920 233
rect 927 226 1144 233
rect 1187 235 1922 237
rect 1177 230 1922 235
rect 1946 239 1962 246
rect 1987 245 2128 252
rect 938 216 960 222
rect 862 207 942 212
rect 1080 206 1185 210
rect 777 195 993 202
rect 1002 195 1058 202
rect 1068 195 1083 202
rect 1092 195 1913 202
rect 780 178 1049 185
rect 1058 178 1128 185
rect 1137 178 1244 185
rect 1107 154 1157 161
rect 1167 155 1385 162
rect 1427 163 1922 165
rect 1417 158 1922 163
rect 1946 167 1962 174
rect 1987 173 2128 180
rect 1374 145 1412 151
rect 1319 134 1428 139
rect 1018 123 1143 130
rect 1152 123 1233 130
rect 1242 123 1298 130
rect 1308 123 1913 130
rect 1020 106 1188 113
rect 1197 106 1289 113
rect 1298 106 1484 113
rect 1353 95 1388 101
rect 1343 82 1398 89
rect 1408 82 1623 89
rect 1667 91 1922 93
rect 1657 86 1922 91
rect 1946 95 1962 102
rect 1987 101 2128 108
rect 1357 69 1676 70
rect 1365 68 1676 69
rect 1365 63 1668 68
rect 1077 51 1323 58
rect 1332 51 1473 58
rect 1482 51 1538 58
rect 1547 51 1920 58
rect 1260 40 1529 41
rect 1260 34 1368 40
rect 1377 34 1529 40
rect 1538 34 1724 41
rect 1473 20 1838 27
rect 1946 23 1962 30
rect 1987 29 2128 36
rect 1586 10 1637 16
rect 1646 10 1866 16
rect -320 -7 -83 0
rect -73 -7 400 0
rect 410 -7 634 0
rect 643 -7 874 0
rect 883 -7 1115 0
rect 1124 -7 1412 0
rect 1421 -7 1607 0
rect 1616 -7 1847 0
rect -320 -18 1335 -11
rect 1341 -12 1567 -11
rect 1341 -18 1402 -12
rect 1408 -18 1567 -12
rect 1574 -18 1650 -11
rect 1658 -18 1920 -11
rect -320 -23 1618 -22
rect -320 -29 1392 -23
rect 1398 -29 1618 -23
rect 1626 -29 1920 -22
rect -320 -34 1590 -33
rect -320 -40 1347 -34
rect 1353 -40 1590 -34
rect 1598 -40 1662 -33
rect 1670 -40 1920 -33
rect -320 -45 1630 -44
rect -320 -51 1381 -45
rect 1387 -51 1630 -45
rect 1638 -51 1920 -44
<< m456contact >>
rect 134 505 149 513
rect 440 434 452 442
rect 646 381 658 390
rect 605 350 620 358
rect 1098 214 1110 222
rect 1141 214 1153 222
rect 1167 214 1179 222
rect 1336 143 1348 151
rect 1335 4 1343 12
<< m6contact >>
rect 136 422 149 430
rect 610 278 618 286
<< metal6 >>
rect 142 430 149 505
rect 142 2 149 422
rect 610 286 617 350
rect 610 1 617 278
rect 651 2 658 381
rect 1102 2 1110 214
rect 1141 2 1149 214
rect 1167 2 1175 214
rect 1341 12 1348 143
rect 1343 4 1348 12
use logic  logic_0
timestamp 1575955143
transform 1 0 -407 0 1 504
box 87 2 327 70
use two_1_mux  two_1_mux_0
timestamp 1575861164
transform 1 0 -125 0 1 565
box 45 -59 125 9
use fadder  fadder_0
timestamp 1575950238
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1575955143
transform 1 0 -87 0 1 432
box 87 2 327 70
use inputff  inputff_0
timestamp 1575939406
transform 1 0 -174 0 1 482
box -76 -120 134 -52
use driver  driver_0
timestamp 1575946641
transform 1 0 -32 0 1 421
box -8 -59 92 9
use fadder  fadder_1
timestamp 1575950238
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1575955143
transform 1 0 153 0 1 360
box 87 2 327 70
use inputff  inputff_1
timestamp 1575939406
transform 1 0 -244 0 1 410
box -76 -120 134 -52
use driver  driver_1
timestamp 1575946641
transform 1 0 -102 0 1 349
box -8 -59 92 9
use inputff  inputff_2
timestamp 1575939406
transform 1 0 66 0 1 410
box -76 -120 134 -52
use driver  driver_2
timestamp 1575946641
transform 1 0 208 0 1 349
box -8 -59 92 9
use fadder  fadder_2
timestamp 1575950238
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1575955143
transform 1 0 393 0 1 288
box 87 2 327 70
use dff  dff_0
timestamp 1575941385
transform 1 0 -320 0 1 279
box 0 -61 150 7
use driver  driver_8
timestamp 1575946641
transform 1 0 -172 0 1 277
box -8 -59 92 9
use inputff  inputff_3
timestamp 1575939406
transform 1 0 -4 0 1 338
box -76 -120 134 -52
use driver  driver_3
timestamp 1575946641
transform 1 0 138 0 1 277
box -8 -59 92 9
use inputff  inputff_4
timestamp 1575939406
transform 1 0 306 0 1 338
box -76 -120 134 -52
use driver  driver_4
timestamp 1575946641
transform 1 0 448 0 1 277
box -8 -59 92 9
use fadder  fadder_3
timestamp 1575950238
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1575955143
transform 1 0 633 0 1 216
box 87 2 327 70
use dff  dff_3
timestamp 1575941385
transform 1 0 -250 0 1 207
box 0 -61 150 7
use driver  driver_11
timestamp 1575946641
transform 1 0 -102 0 1 205
box -8 -59 92 9
use dff  dff_2
timestamp 1575941385
transform 1 0 -10 0 1 207
box 0 -61 150 7
use driver  driver_10
timestamp 1575946641
transform 1 0 138 0 1 205
box -8 -59 92 9
use dff  dff_1
timestamp 1575941385
transform 1 0 230 0 1 207
box 0 -61 150 7
use driver  driver_9
timestamp 1575946641
transform 1 0 378 0 1 205
box -8 -59 92 9
use inputff  inputff_5
timestamp 1575939406
transform 1 0 546 0 1 266
box -76 -120 134 -52
use driver  driver_5
timestamp 1575946641
transform 1 0 688 0 1 205
box -8 -59 92 9
use fadder  fadder_4
timestamp 1575950238
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1575955143
transform 1 0 873 0 1 144
box 87 2 327 70
use inputff  inputff_6
timestamp 1575939406
transform 1 0 786 0 1 194
box -76 -120 134 -52
use driver  driver_6
timestamp 1575946641
transform 1 0 928 0 1 133
box -8 -59 92 9
use fadder  fadder_5
timestamp 1575950238
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1575955143
transform 1 0 1113 0 1 72
box 87 2 327 70
use inputff  inputff_7
timestamp 1575939406
transform 1 0 846 0 1 122
box -76 -120 134 -52
use driver  driver_7
timestamp 1575946641
transform 1 0 988 0 1 61
box -8 -59 92 9
use fadder  fadder_6
timestamp 1575950238
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1575950238
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1575955143
transform 1 0 1353 0 1 0
box 87 2 327 70
use inv_9_6  inv_9_6_0
array 0 0 30 0 7 72
timestamp 1575941223
transform 1 0 1920 0 1 62
box 0 -60 30 8
use enff  enff_0
array 0 0 191 0 7 72
timestamp 1575941385
transform 1 0 1993 0 1 2
box -43 0 147 68
use mult  mult_0
timestamp 1575939595
transform 1 0 241 0 1 432
box -241 -432 1689 142
<< labels >>
rlabel m4contact 430 469 430 469 1 4mux_to_2mux_1
rlabel metal5 -318 558 -318 558 3 y0
rlabel metal5 -177 486 -177 486 1 y1
rlabel metal5 63 414 63 414 1 y2
rlabel metal5 304 342 304 342 1 y3
rlabel metal5 544 271 544 271 1 y4
rlabel metal5 784 199 784 199 1 y5
rlabel metal5 1025 126 1025 126 1 y6
rlabel metal5 1084 55 1084 55 1 y7
rlabel metal5 -317 -3 -317 -3 3 opcode2
rlabel m4contact -8 535 -8 535 1 nz0
rlabel metal5 1659 88 1659 88 1 nz6
rlabel metal3 1918 25 1918 25 1 nz7
rlabel m345contact 459 448 459 448 1 nz1
rlabel m345contact 700 380 700 380 1 nz2
rlabel m345contact 941 308 941 308 1 nz3
rlabel metal5 1181 233 1181 233 1 nz4
rlabel metal5 1420 160 1420 160 1 nz5
rlabel metal5 2123 537 2123 537 1 z0
rlabel metal5 2123 465 2123 465 1 z1
rlabel metal5 2123 392 2123 392 1 z2
rlabel metal5 2123 321 2123 321 1 z3
rlabel metal5 2123 248 2123 248 1 z4
rlabel metal5 2123 176 2123 176 1 z5
rlabel metal5 2123 105 2123 105 1 z6
rlabel metal5 2123 32 2123 32 1 z7
rlabel metal4 1954 546 1954 546 1 c_en
rlabel m2contact 2189 510 2189 510 1 Gnd
rlabel metal1 2210 511 2210 511 7 Vdd
rlabel m5contact 1824 582 1824 582 1 clk
rlabel metal4 239 580 239 580 1 x0
rlabel metal4 1439 580 1439 580 1 x5
rlabel metal4 1679 581 1679 581 1 x6
rlabel metal4 1920 581 1920 581 1 x7
rlabel metal4 1199 581 1199 581 1 x4
rlabel metal4 959 580 959 580 1 x3
rlabel metal4 718 590 718 590 1 x2
rlabel metal4 479 576 479 576 1 x1
rlabel metal3 -318 251 -318 251 3 Actrl
rlabel metal4 233 -39 233 -39 1 opcode2
rlabel metal5 1639 -26 1639 -26 1 opcode0
rlabel metal5 1639 -37 1639 -37 1 opcode1n
rlabel metal5 1639 -48 1639 -48 1 opcode0n
rlabel metal5 1639 -15 1639 -15 1 opcode1
<< end >>
