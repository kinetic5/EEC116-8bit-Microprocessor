magic
tech scmos
timestamp 1576013433
<< ntransistor >>
rect 14 -38 16 -34
rect 24 -38 26 -34
rect 34 -38 36 -34
rect 44 -38 46 -34
rect 64 -38 66 -34
rect 74 -38 76 -34
rect 84 -38 86 -34
rect 94 -38 96 -34
rect 54 -46 56 -42
rect 114 -38 116 -34
rect 104 -46 106 -42
rect 124 -42 126 -34
rect 134 -42 136 -34
<< ptransistor >>
rect 54 -12 56 -6
rect 14 -22 16 -16
rect 24 -22 26 -16
rect 34 -22 36 -16
rect 44 -22 46 -16
rect 104 -12 106 -6
rect 64 -22 66 -16
rect 74 -22 76 -16
rect 84 -22 86 -16
rect 94 -22 96 -16
rect 114 -22 116 -16
rect 124 -22 126 -10
rect 134 -22 136 -10
<< ndiffusion >>
rect 13 -38 14 -34
rect 16 -38 17 -34
rect 23 -38 24 -34
rect 26 -38 27 -34
rect 33 -38 34 -34
rect 36 -38 37 -34
rect 43 -38 44 -34
rect 46 -38 47 -34
rect 63 -38 64 -34
rect 66 -38 67 -34
rect 73 -38 74 -34
rect 76 -38 77 -34
rect 83 -38 84 -34
rect 86 -38 87 -34
rect 93 -38 94 -34
rect 96 -38 97 -34
rect 57 -42 62 -38
rect 49 -46 54 -42
rect 56 -46 62 -42
rect 49 -50 53 -46
rect 113 -38 114 -34
rect 116 -38 124 -34
rect 99 -46 104 -42
rect 106 -46 107 -42
rect 99 -50 103 -46
rect 117 -42 124 -38
rect 126 -35 134 -34
rect 126 -42 127 -35
rect 133 -42 134 -35
rect 136 -42 137 -34
rect 117 -43 123 -42
<< pdiffusion >>
rect 53 -12 54 -6
rect 56 -12 62 -6
rect 13 -22 14 -16
rect 16 -22 17 -16
rect 23 -22 24 -16
rect 26 -22 27 -16
rect 33 -22 34 -16
rect 36 -22 37 -16
rect 43 -22 44 -16
rect 46 -22 47 -16
rect 57 -16 62 -12
rect 103 -12 104 -6
rect 106 -11 107 -6
rect 106 -12 113 -11
rect 63 -22 64 -16
rect 66 -22 67 -16
rect 73 -22 74 -16
rect 76 -22 77 -16
rect 83 -22 84 -16
rect 86 -22 87 -16
rect 93 -22 94 -16
rect 96 -22 97 -16
rect 123 -13 124 -10
rect 117 -16 124 -13
rect 113 -22 114 -16
rect 116 -22 124 -16
rect 126 -21 127 -10
rect 133 -21 134 -10
rect 126 -22 134 -21
rect 136 -22 137 -10
<< ndcontact >>
rect 7 -38 13 -34
rect 17 -38 23 -34
rect 27 -38 33 -34
rect 37 -38 43 -34
rect 47 -38 53 -34
rect 57 -38 63 -34
rect 67 -38 73 -34
rect 77 -38 83 -34
rect 87 -38 93 -34
rect 97 -38 102 -34
rect 107 -38 113 -34
rect 137 -42 143 -34
rect 117 -48 123 -43
rect 49 -54 53 -50
rect 99 -54 103 -50
<< pdcontact >>
rect 47 -12 53 -6
rect 7 -22 13 -16
rect 17 -22 23 -16
rect 27 -22 33 -16
rect 37 -22 43 -16
rect 47 -22 53 -16
rect 97 -12 103 -6
rect 57 -22 63 -16
rect 67 -22 73 -16
rect 77 -22 83 -16
rect 87 -22 93 -16
rect 97 -22 102 -16
rect 117 -13 123 -8
rect 107 -22 113 -16
rect 137 -22 143 -10
<< polysilicon >>
rect 4 -50 6 -4
rect 14 -6 16 -4
rect 24 -6 26 -4
rect 14 -16 16 -12
rect 24 -16 26 -12
rect 34 -16 36 -4
rect 44 -16 46 -4
rect 54 -6 56 -3
rect 64 -6 66 -4
rect 74 -6 76 -4
rect 14 -25 16 -22
rect 24 -25 26 -22
rect 34 -25 36 -22
rect 14 -34 16 -31
rect 24 -34 26 -31
rect 34 -34 36 -31
rect 44 -34 46 -22
rect 54 -25 56 -12
rect 64 -16 66 -12
rect 74 -16 76 -12
rect 84 -16 86 -4
rect 94 -16 96 -4
rect 104 -6 106 -3
rect 64 -25 66 -22
rect 74 -25 76 -22
rect 84 -25 86 -22
rect 14 -42 16 -38
rect 24 -42 26 -38
rect 14 -50 16 -48
rect 24 -50 26 -48
rect 34 -50 36 -38
rect 44 -41 46 -38
rect 54 -42 56 -31
rect 64 -34 66 -31
rect 74 -34 76 -31
rect 84 -34 86 -31
rect 94 -34 96 -22
rect 104 -25 106 -12
rect 114 -16 116 -4
rect 124 -10 126 -4
rect 134 -10 136 -4
rect 114 -25 116 -22
rect 124 -25 126 -22
rect 134 -25 136 -22
rect 64 -42 66 -38
rect 74 -42 76 -38
rect 44 -50 46 -46
rect 54 -50 56 -46
rect 64 -50 66 -48
rect 74 -49 76 -48
rect 84 -49 86 -38
rect 94 -41 96 -38
rect 104 -42 106 -31
rect 114 -34 116 -31
rect 124 -34 126 -31
rect 134 -34 136 -31
rect 94 -49 96 -46
rect 104 -49 106 -46
rect 114 -49 116 -38
rect 124 -49 126 -42
rect 134 -50 136 -42
rect 144 -50 146 -4
<< polycontact >>
rect 34 -31 38 -25
rect 52 -31 56 -25
rect 84 -31 88 -25
rect 104 -31 108 -25
rect 122 -31 127 -25
rect 133 -31 138 -25
<< metal1 >>
rect 0 -1 150 7
rect 37 -16 43 -1
rect 47 -6 53 -1
rect 87 -16 93 -1
rect 97 -6 103 -1
rect 117 -8 123 -1
rect 137 -10 143 -1
rect 7 -24 13 -22
rect 7 -34 13 -32
rect 17 -29 23 -22
rect 26 -22 27 -16
rect 26 -34 31 -22
rect 47 -25 53 -22
rect 38 -31 52 -25
rect 47 -34 53 -31
rect 59 -34 63 -22
rect 26 -38 27 -34
rect 36 -38 37 -34
rect 67 -27 73 -22
rect 67 -34 73 -32
rect 76 -22 77 -16
rect 105 -22 107 -16
rect 113 -21 117 -16
rect 113 -22 123 -21
rect 76 -34 81 -22
rect 97 -25 101 -22
rect 105 -25 109 -22
rect 88 -31 94 -25
rect 108 -31 109 -25
rect 97 -34 101 -31
rect 105 -34 109 -31
rect 76 -38 77 -34
rect 86 -38 87 -34
rect 105 -38 107 -34
rect 113 -35 123 -34
rect 113 -38 117 -35
rect 36 -53 40 -38
rect 0 -54 49 -53
rect 86 -53 90 -38
rect 105 -39 117 -38
rect 53 -54 99 -53
rect 117 -53 123 -48
rect 137 -53 143 -42
rect 103 -54 150 -53
rect 0 -61 150 -54
<< pm12contact >>
rect 13 -12 18 -6
rect 22 -12 27 -6
rect 63 -12 68 -6
rect 72 -12 77 -6
rect 112 -31 118 -25
rect 13 -48 18 -42
rect 22 -48 27 -42
rect 43 -46 48 -41
rect 63 -48 68 -42
rect 72 -48 77 -42
rect 93 -46 98 -41
<< pdm12contact >>
rect 107 -11 113 -6
rect 127 -21 133 -10
<< ndm12contact >>
rect 127 -42 133 -35
rect 107 -47 113 -42
<< metal2 >>
rect 12 -2 113 4
rect 12 -6 18 -2
rect 72 -6 78 -2
rect 12 -12 13 -6
rect 77 -12 78 -6
rect 83 -6 113 -2
rect 43 -41 48 -39
rect 27 -48 28 -42
rect 22 -52 28 -48
rect 62 -48 63 -42
rect 62 -52 68 -48
rect 83 -52 89 -6
rect 103 -21 112 -15
rect 106 -31 112 -21
rect 93 -41 98 -40
rect 107 -52 113 -47
rect 13 -58 113 -52
<< m3contact >>
rect 27 -12 33 -6
rect 57 -12 63 -6
rect 43 -39 48 -34
rect 7 -48 13 -42
rect 72 -42 78 -37
rect 127 -10 133 -3
rect 95 -21 103 -13
rect 93 -40 98 -35
rect 127 -49 133 -42
<< m123contact >>
rect 7 -32 13 -24
rect 17 -34 23 -29
rect 67 -32 73 -27
rect 117 -21 123 -16
rect 94 -31 101 -25
rect 127 -31 133 -25
rect 117 -40 123 -35
<< metal3 >>
rect 27 -2 123 4
rect 27 -6 33 -2
rect 57 -6 63 -2
rect 117 -16 123 -2
rect 133 -10 143 -3
rect 67 -27 90 -24
rect 73 -29 90 -27
rect 17 -38 43 -34
rect 85 -35 90 -29
rect 101 -31 127 -25
rect 85 -39 93 -35
rect 87 -40 93 -39
rect 72 -44 78 -42
rect 117 -44 123 -40
rect 137 -42 143 -10
rect 13 -48 123 -44
rect 7 -49 123 -48
rect 133 -49 143 -42
<< labels >>
rlabel metal3 141 -28 141 -28 1 q
rlabel m123contact 10 -28 10 -28 1 d
rlabel m123contact 70 -29 70 -29 1 transm23_out
rlabel metal1 20 -27 20 -27 1 transm01_out
rlabel pdm12contact 110 -9 110 -9 1 _clk
rlabel m3contact 99 -14 99 -14 1 clk
rlabel metal1 5 3 5 3 4 Vdd
rlabel metal1 4 -56 4 -56 2 Gnd
rlabel metal1 107 -33 107 -33 1 _nclk
<< end >>
