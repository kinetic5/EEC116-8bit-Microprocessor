magic
tech scmos
timestamp 1575856977
<< error_s >>
rect -217 540 -211 546
rect -148 536 -142 538
rect 23 468 29 474
rect 92 464 98 466
rect 263 396 269 402
rect 503 324 509 330
rect 743 252 749 258
rect 983 180 989 186
rect 1223 108 1229 114
rect 1463 36 1469 42
<< metal2 >>
rect -13 441 -7 455
rect -13 435 73 441
rect 67 427 73 435
rect 227 369 233 383
rect 227 363 313 369
rect 307 349 313 363
rect 467 297 473 313
rect 467 291 553 297
rect 547 278 553 291
rect 707 225 713 239
rect 707 219 793 225
rect 787 206 793 219
rect 947 153 953 168
rect 947 147 1033 153
rect 1027 133 1033 147
rect 1187 69 1193 95
rect 1147 63 1193 69
rect 1247 61 1273 67
rect 1247 44 1253 61
<< m3contact >>
rect -173 543 -167 549
rect 67 471 73 477
rect 307 399 313 405
rect 547 327 553 333
rect 787 255 793 261
rect 1027 183 1033 189
rect 1267 111 1273 117
rect 1507 39 1513 45
<< metal3 >>
rect -163 553 -141 557
rect 0 558 8 563
rect -207 546 -201 553
rect -163 551 -132 553
rect -167 543 -151 544
rect -173 538 -151 543
rect -138 538 -132 551
rect 2 510 8 558
rect 12 538 18 552
rect 252 538 258 552
rect 492 538 498 552
rect 732 538 738 552
rect 972 538 978 552
rect 1212 538 1218 552
rect 1452 538 1458 552
rect 1692 538 1698 552
rect -3 501 3 510
rect -83 495 3 501
rect -83 477 -77 495
rect 83 481 99 485
rect 239 486 247 491
rect 33 474 39 481
rect 83 479 108 481
rect 73 471 89 472
rect 67 466 89 471
rect 102 463 108 479
rect 242 438 247 486
rect 237 432 247 438
rect 237 429 243 432
rect 157 423 243 429
rect 157 406 163 423
rect 323 409 339 413
rect 479 414 487 419
rect 273 402 279 409
rect 323 407 348 409
rect 313 399 329 400
rect 307 394 329 399
rect 342 391 348 407
rect 482 366 487 414
rect 476 360 488 366
rect 476 357 482 360
rect 387 351 482 357
rect 387 333 393 351
rect 563 337 579 341
rect 718 342 727 347
rect 513 330 519 337
rect 563 335 588 337
rect 553 327 569 328
rect 547 322 569 327
rect 582 319 588 335
rect 722 294 727 342
rect 717 288 728 294
rect 717 285 723 288
rect 637 279 723 285
rect 637 261 643 279
rect 803 265 819 269
rect 952 270 967 275
rect 753 258 759 265
rect 803 263 828 265
rect 793 255 809 256
rect 787 250 809 255
rect 822 247 828 263
rect 962 222 967 270
rect 957 216 968 222
rect 957 213 963 216
rect 877 207 963 213
rect 877 190 883 207
rect 1043 193 1059 197
rect 1192 198 1207 203
rect 993 186 999 193
rect 1043 191 1068 193
rect 1033 183 1049 184
rect 1027 178 1049 183
rect 1062 173 1068 191
rect 1202 150 1207 198
rect 1196 144 1208 150
rect 1196 141 1202 144
rect 1117 135 1202 141
rect 1117 118 1123 135
rect 1283 121 1299 125
rect 1428 126 1436 134
rect 1233 114 1239 121
rect 1283 119 1308 121
rect 1273 111 1289 112
rect 1267 106 1289 111
rect 1302 101 1308 119
rect 1177 45 1183 62
rect 1357 45 1363 63
rect 1523 49 1539 53
rect 1668 54 1676 62
rect 1473 42 1479 49
rect 1523 47 1548 49
rect 1513 39 1529 40
rect 1507 34 1529 39
rect 1542 34 1548 47
<< m4contact >>
rect 286 533 296 543
rect 526 533 536 543
rect 766 533 776 543
rect 1006 533 1016 543
rect 1246 533 1256 543
rect 1486 533 1496 543
rect 1726 533 1736 543
rect -117 463 -108 472
rect -72 463 -63 472
rect 123 391 132 400
rect 168 391 177 400
rect 363 319 372 328
rect 408 319 417 328
rect 603 246 612 255
rect 648 247 657 256
rect 843 174 852 183
rect 888 175 897 184
rect 1083 103 1092 112
rect 1128 103 1137 112
rect 1177 62 1185 68
rect 1143 31 1152 40
rect 1188 31 1197 40
rect 1323 31 1332 40
<< metal4 >>
rect -115 472 -108 553
rect -70 472 -63 536
rect 125 400 132 481
rect 289 475 296 533
rect 170 400 177 464
rect 365 328 372 409
rect 529 403 536 533
rect 410 328 417 392
rect 605 255 612 337
rect 769 331 776 533
rect 650 256 657 320
rect 845 183 852 265
rect 1009 259 1016 533
rect 890 184 897 248
rect 1085 112 1092 193
rect 1249 187 1256 533
rect 1130 112 1137 176
rect 1145 40 1152 121
rect 1177 68 1184 134
rect 1489 115 1496 533
rect 1190 40 1197 104
rect 1323 40 1332 49
rect 1729 43 1736 533
<< m345contact >>
rect -207 553 -198 562
rect -141 553 -132 562
rect -220 538 -211 547
rect -151 536 -142 545
rect 12 552 22 562
rect 252 552 262 562
rect 492 552 502 562
rect 732 552 742 562
rect 972 552 982 562
rect 1212 552 1222 562
rect 1452 552 1462 562
rect 1692 552 1702 562
rect 46 533 56 543
rect 33 481 42 490
rect 99 481 108 490
rect 20 466 29 475
rect 89 464 98 473
rect 273 409 282 418
rect 339 409 348 418
rect 260 394 269 403
rect 329 394 338 403
rect 513 337 522 346
rect 579 337 588 346
rect 500 322 509 331
rect 569 322 578 331
rect 753 265 762 274
rect 819 265 828 274
rect 740 250 749 259
rect 809 250 818 259
rect 993 193 1002 202
rect 1059 193 1068 202
rect 980 178 989 187
rect 1049 178 1058 187
rect 1428 134 1436 140
rect 1233 121 1242 130
rect 1299 121 1308 130
rect 1220 106 1229 115
rect 1289 106 1298 115
rect 1357 63 1365 69
rect 1668 62 1676 68
rect 1473 49 1482 58
rect 1539 49 1548 58
rect 1368 31 1377 40
rect 1460 34 1469 43
rect 1529 34 1538 43
<< m5contact >>
rect -117 553 -108 562
rect -72 536 -63 545
rect 123 481 132 490
rect 168 464 177 473
rect 287 466 296 475
rect 363 409 372 418
rect 408 392 417 401
rect 527 394 536 403
rect 603 337 612 346
rect 648 320 657 329
rect 767 322 776 331
rect 843 265 852 274
rect 888 248 897 257
rect 1007 250 1016 259
rect 1083 193 1092 202
rect 1128 176 1137 185
rect 1247 178 1256 187
rect 1177 134 1185 140
rect 1143 121 1152 130
rect 1188 104 1197 113
rect 1487 106 1496 115
rect 1323 49 1332 58
rect 1727 34 1736 43
<< metal5 >>
rect -240 555 -207 562
rect -198 555 -141 562
rect -132 555 -117 562
rect -108 555 12 562
rect 22 555 252 562
rect 262 555 492 562
rect 502 555 732 562
rect 742 555 972 562
rect 982 555 1212 562
rect 1222 555 1452 562
rect 1462 555 1692 562
rect 1702 555 1913 562
rect -240 538 -220 545
rect -211 538 -151 545
rect -142 538 -72 545
rect -63 543 56 545
rect -63 538 46 543
rect -180 483 0 490
rect 1 483 33 490
rect 42 483 99 490
rect 108 483 123 490
rect 132 483 1920 490
rect -180 466 20 473
rect 29 466 89 473
rect 98 466 168 473
rect 177 466 287 473
rect 60 411 273 418
rect 282 411 339 418
rect 348 411 363 418
rect 372 411 1913 418
rect 60 394 260 401
rect 269 394 329 401
rect 338 394 408 401
rect 417 394 527 401
rect 300 339 513 346
rect 522 339 579 346
rect 588 339 603 346
rect 612 339 1913 346
rect 300 322 500 329
rect 509 322 569 329
rect 578 322 648 329
rect 657 322 767 329
rect 540 267 753 274
rect 762 267 819 274
rect 828 267 843 274
rect 852 267 1913 274
rect 540 250 740 257
rect 749 250 809 257
rect 818 250 888 257
rect 897 250 1007 257
rect 780 195 993 202
rect 1002 195 1059 202
rect 1068 195 1083 202
rect 1092 195 1913 202
rect 780 178 980 185
rect 989 178 1049 185
rect 1058 178 1128 185
rect 1137 178 1247 185
rect 1177 140 1436 141
rect 1185 134 1428 140
rect 1020 123 1143 130
rect 1152 123 1233 130
rect 1242 123 1299 130
rect 1308 123 1913 130
rect 1020 106 1188 113
rect 1197 106 1220 113
rect 1229 106 1289 113
rect 1298 106 1487 113
rect 1357 69 1676 70
rect 1365 68 1676 69
rect 1365 63 1668 68
rect 1080 51 1323 58
rect 1332 51 1440 58
rect 1442 51 1473 58
rect 1482 51 1539 58
rect 1548 51 1920 58
rect 1260 40 1460 41
rect 1260 34 1368 40
rect 1377 34 1460 40
rect 1469 34 1529 41
rect 1538 34 1727 41
<< metal6 >>
rect 1874 62 1882 593
rect 1890 2 1898 593
use logic  logic_0
timestamp 1575855885
transform 1 0 -327 0 1 504
box 87 2 327 70
use fadder  fadder_0
timestamp 1575778664
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1575855885
transform 1 0 -87 0 1 432
box 87 2 327 70
use fadder  fadder_1
timestamp 1575778664
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1575855885
transform 1 0 153 0 1 360
box 87 2 327 70
use fadder  fadder_2
timestamp 1575778664
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1575855885
transform 1 0 393 0 1 288
box 87 2 327 70
use fadder  fadder_3
timestamp 1575778664
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1575855885
transform 1 0 633 0 1 216
box 87 2 327 70
use fadder  fadder_4
timestamp 1575778664
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1575855885
transform 1 0 873 0 1 144
box 87 2 327 70
use fadder  fadder_5
timestamp 1575778664
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1575855885
transform 1 0 1113 0 1 72
box 87 2 327 70
use fadder  fadder_6
timestamp 1575778664
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1575778664
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1575855885
transform 1 0 1353 0 1 0
box 87 2 327 70
use mult  mult_0
timestamp 1575856188
transform 1 0 241 0 1 432
box -241 -432 1679 142
<< labels >>
rlabel metal6 1878 590 1878 590 5 Vdd
rlabel metal6 1894 589 1894 589 5 Gnd
<< end >>
