magic
tech scmos
timestamp 1576123792
<< error_p >>
rect 17 34 23 35
rect 37 34 43 35
rect 57 34 63 35
rect 67 34 113 35
<< nwell >>
rect 0 52 230 102
<< pwell >>
rect 0 -2 230 40
<< ntransistor >>
rect 14 27 16 33
rect 24 27 26 33
rect 34 24 36 33
rect 44 24 46 33
rect 54 24 56 33
rect 64 24 66 33
rect 74 20 76 35
rect 84 20 86 35
rect 94 20 96 35
rect 104 20 106 35
rect 124 17 126 34
rect 134 17 136 34
rect 144 17 146 34
rect 154 17 156 34
rect 164 17 166 34
rect 174 17 176 34
rect 184 17 186 34
rect 194 17 196 34
rect 204 17 206 34
rect 214 17 216 34
<< ptransistor >>
rect 14 68 16 80
rect 24 68 26 80
rect 34 66 36 80
rect 44 66 46 80
rect 54 66 56 80
rect 64 66 66 80
rect 74 61 76 84
rect 84 61 86 84
rect 94 61 96 84
rect 104 61 106 84
rect 124 58 126 83
rect 134 58 136 83
rect 144 58 146 83
rect 154 58 156 83
rect 164 58 166 83
rect 174 58 176 83
rect 184 58 186 83
rect 194 58 196 83
rect 204 58 206 83
rect 214 58 216 83
<< ndiffusion >>
rect 13 27 14 33
rect 16 27 17 33
rect 23 27 24 33
rect 26 27 27 33
rect 33 24 34 33
rect 36 24 37 33
rect 43 24 44 33
rect 46 24 47 33
rect 53 24 54 33
rect 56 24 57 33
rect 63 24 64 33
rect 66 24 67 33
rect 73 20 74 35
rect 76 20 77 35
rect 83 20 84 35
rect 86 20 87 35
rect 93 20 94 35
rect 96 20 97 35
rect 103 20 104 35
rect 106 20 107 35
rect 123 17 124 34
rect 126 17 127 34
rect 133 17 134 34
rect 136 17 137 34
rect 143 17 144 34
rect 146 17 147 34
rect 153 17 154 34
rect 156 17 157 34
rect 163 17 164 34
rect 166 17 167 34
rect 173 17 174 34
rect 176 17 177 34
rect 183 17 184 34
rect 186 17 187 34
rect 193 17 194 34
rect 196 17 197 34
rect 203 17 204 34
rect 206 17 207 34
rect 213 17 214 34
rect 216 17 217 34
<< pdiffusion >>
rect 13 68 14 80
rect 16 68 17 80
rect 23 68 24 80
rect 26 68 27 80
rect 33 66 34 80
rect 36 66 37 80
rect 43 66 44 80
rect 46 66 47 80
rect 53 66 54 80
rect 56 66 57 80
rect 63 66 64 80
rect 66 66 67 80
rect 73 61 74 84
rect 76 62 77 84
rect 83 62 84 84
rect 76 61 84 62
rect 86 61 87 84
rect 93 61 94 84
rect 96 62 97 84
rect 103 62 104 84
rect 96 61 104 62
rect 106 61 107 84
rect 123 58 124 83
rect 126 58 127 83
rect 133 58 134 83
rect 136 58 137 83
rect 143 58 144 83
rect 146 58 147 83
rect 153 58 154 83
rect 156 58 157 83
rect 163 58 164 83
rect 166 58 167 83
rect 173 58 174 83
rect 176 58 177 83
rect 183 58 184 83
rect 186 58 187 83
rect 193 58 194 83
rect 196 58 197 83
rect 203 58 204 83
rect 206 58 207 83
rect 213 58 214 83
rect 216 58 217 83
<< ndcontact >>
rect 7 25 13 33
rect 27 24 33 33
rect 47 24 53 33
rect 67 20 73 35
rect 87 20 93 35
rect 107 20 113 35
rect 117 17 123 34
rect 137 17 143 34
rect 157 17 163 34
rect 177 17 183 34
rect 197 17 203 34
rect 217 17 223 34
<< pdcontact >>
rect 7 68 13 80
rect 27 66 33 80
rect 47 66 53 80
rect 67 61 73 84
rect 87 61 93 84
rect 107 61 113 84
rect 117 58 123 83
rect 137 58 143 83
rect 157 58 163 83
rect 177 58 183 83
rect 197 58 203 83
rect 217 58 223 83
<< polysilicon >>
rect 4 14 6 86
rect 14 80 16 86
rect 24 80 26 86
rect 34 80 36 86
rect 44 80 46 86
rect 54 80 56 86
rect 64 80 66 86
rect 74 84 76 87
rect 84 84 86 87
rect 94 84 96 87
rect 104 84 106 87
rect 14 58 16 68
rect 24 58 26 68
rect 34 58 36 66
rect 44 58 46 66
rect 54 58 56 66
rect 64 58 66 66
rect 74 58 76 61
rect 84 58 86 61
rect 94 58 96 61
rect 104 58 106 61
rect 12 45 13 58
rect 14 33 16 45
rect 14 14 16 27
rect 24 33 26 45
rect 34 33 36 45
rect 24 14 26 27
rect 44 33 46 45
rect 54 33 56 45
rect 34 14 36 22
rect 44 14 46 22
rect 64 33 66 45
rect 74 35 76 45
rect 84 35 86 45
rect 94 35 96 45
rect 104 35 106 45
rect 54 14 56 22
rect 64 14 66 22
rect 74 14 76 20
rect 84 14 86 20
rect 94 14 96 20
rect 104 14 106 20
rect 114 14 116 86
rect 124 83 126 86
rect 134 83 136 86
rect 144 83 146 86
rect 154 83 156 86
rect 164 83 166 86
rect 174 83 176 86
rect 184 83 186 86
rect 194 83 196 86
rect 204 83 206 86
rect 214 83 216 86
rect 124 54 126 58
rect 134 54 136 58
rect 144 54 146 58
rect 154 54 156 58
rect 164 54 166 58
rect 174 54 176 58
rect 184 54 186 58
rect 194 54 196 58
rect 204 54 206 58
rect 214 54 216 58
rect 124 34 126 38
rect 134 34 136 38
rect 144 34 146 38
rect 154 34 156 38
rect 164 34 166 38
rect 174 34 176 38
rect 184 34 186 38
rect 194 34 196 38
rect 204 34 206 38
rect 214 34 216 38
rect 124 14 126 17
rect 134 14 136 17
rect 144 14 146 17
rect 154 14 156 17
rect 164 14 166 17
rect 174 14 176 17
rect 184 14 186 17
rect 194 14 196 17
rect 204 14 206 17
rect 214 14 216 17
rect 224 14 226 86
<< polycontact >>
rect 13 45 18 58
rect 22 45 28 58
rect 42 45 48 58
rect 52 45 58 58
rect 62 45 68 58
rect 82 45 88 58
rect 92 45 98 58
rect 102 45 108 58
rect 132 38 138 54
rect 142 38 148 54
rect 152 38 158 54
rect 162 38 168 54
rect 172 38 178 54
rect 182 38 188 54
rect 192 38 198 54
rect 202 38 208 54
rect 212 38 218 54
<< polynplus >>
rect 34 22 36 24
rect 44 22 46 24
rect 54 22 56 24
rect 64 22 66 24
<< metal1 >>
rect 0 88 230 100
rect 7 80 13 88
rect 27 80 33 88
rect 47 80 53 88
rect 67 84 73 88
rect 87 84 93 88
rect 107 84 113 88
rect 117 83 123 88
rect 137 83 143 88
rect 157 83 163 88
rect 177 83 183 88
rect 197 83 203 88
rect 217 83 223 88
rect 18 45 22 58
rect 38 45 42 58
rect 48 45 52 58
rect 58 45 62 58
rect 78 45 82 58
rect 88 45 92 58
rect 98 45 102 58
rect 128 38 132 54
rect 138 38 142 54
rect 148 38 152 54
rect 158 38 162 54
rect 168 38 172 54
rect 178 38 182 54
rect 188 38 192 54
rect 198 38 202 54
rect 208 38 212 54
rect 7 12 13 25
rect 27 12 33 24
rect 47 12 53 24
rect 67 12 73 20
rect 87 12 93 20
rect 107 12 113 20
rect 117 12 123 17
rect 137 12 143 17
rect 157 12 163 17
rect 177 12 183 17
rect 197 12 203 17
rect 217 12 223 17
rect 0 0 230 12
<< pm12contact >>
rect 32 45 38 58
rect 72 45 78 58
rect 122 38 128 54
<< pdm12contact >>
rect 17 68 23 80
rect 37 66 43 80
rect 57 66 63 80
rect 77 62 83 84
rect 97 62 103 84
rect 127 58 133 83
rect 147 58 153 83
rect 167 58 173 83
rect 187 58 193 83
rect 207 58 213 83
<< ndm12contact >>
rect 17 23 23 35
rect 37 23 43 35
rect 57 23 63 35
rect 77 20 83 35
rect 97 20 103 35
rect 127 17 133 34
rect 147 17 153 34
rect 167 17 173 34
rect 187 17 193 34
rect 207 17 213 34
<< metal2 >>
rect 23 68 25 80
rect 17 58 25 68
rect 43 66 57 80
rect 49 58 63 66
rect 83 62 97 84
rect 103 62 107 84
rect 17 45 32 58
rect 49 45 72 58
rect 93 54 107 62
rect 133 58 147 83
rect 153 58 167 83
rect 173 58 187 83
rect 193 58 207 83
rect 17 35 25 45
rect 49 35 63 45
rect 93 38 122 54
rect 93 35 107 38
rect 23 23 25 35
rect 43 23 57 35
rect 83 20 97 35
rect 103 20 107 35
rect 190 34 214 58
rect 133 17 147 34
rect 153 17 167 34
rect 173 17 187 34
rect 193 17 207 34
<< m3contact >>
rect 214 34 228 58
<< m123contact >>
rect 4 40 13 63
<< labels >>
rlabel m123contact 8 51 8 51 1 in
rlabel m3contact 227 45 227 45 7 out
rlabel metal1 75 92 75 92 1 Vdd
rlabel metal1 73 3 73 3 1 Gnd
<< end >>
