magic
tech scmos
timestamp 1576133447
<< nwell >>
rect 6 42 257 79
rect 6 40 175 42
<< pwell >>
rect 175 40 245 42
rect 6 7 246 40
<< ntransistor >>
rect 20 30 22 34
rect 30 30 32 34
rect 50 28 52 34
rect 60 25 62 34
rect 70 28 72 34
rect 80 28 82 34
rect 100 28 102 34
rect 120 28 122 34
rect 130 28 132 34
rect 150 25 152 34
rect 190 30 192 36
rect 200 32 202 36
rect 180 21 182 25
rect 220 28 222 36
rect 230 28 232 36
<< ptransistor >>
rect 20 46 22 52
rect 30 46 32 52
rect 50 46 52 55
rect 60 46 62 58
rect 70 46 72 55
rect 80 46 82 55
rect 100 46 102 55
rect 120 46 122 52
rect 130 46 132 52
rect 150 46 152 58
rect 180 59 182 65
rect 190 48 192 54
rect 200 48 202 54
rect 220 48 222 60
rect 230 48 232 60
<< ndiffusion >>
rect 19 30 20 34
rect 22 30 30 34
rect 32 33 39 34
rect 32 30 33 33
rect 43 33 50 34
rect 49 28 50 33
rect 52 28 53 34
rect 59 25 60 34
rect 62 28 63 34
rect 69 28 70 34
rect 72 29 73 34
rect 79 29 80 34
rect 72 28 80 29
rect 82 28 83 34
rect 62 25 66 28
rect 99 28 100 34
rect 102 28 103 34
rect 119 28 120 34
rect 122 28 130 34
rect 132 33 139 34
rect 132 28 133 33
rect 149 25 150 34
rect 152 25 153 34
rect 183 34 190 36
rect 183 30 184 34
rect 189 30 190 34
rect 192 32 194 36
rect 199 32 200 36
rect 202 32 203 36
rect 192 30 196 32
rect 178 24 180 25
rect 173 21 180 24
rect 182 21 188 25
rect 183 17 188 21
rect 219 29 220 36
rect 213 28 220 29
rect 222 28 223 36
rect 229 28 230 36
rect 232 28 233 36
<< pdiffusion >>
rect 19 46 20 52
rect 22 47 23 52
rect 29 47 30 52
rect 22 46 30 47
rect 32 46 33 52
rect 49 47 50 55
rect 43 46 50 47
rect 52 46 53 55
rect 59 46 60 58
rect 62 55 66 58
rect 62 46 63 55
rect 69 46 70 55
rect 72 52 80 55
rect 72 46 73 52
rect 79 46 80 52
rect 82 52 86 55
rect 82 46 83 52
rect 93 54 100 55
rect 99 46 100 54
rect 102 46 103 55
rect 119 46 120 52
rect 122 47 123 52
rect 129 47 130 52
rect 122 46 130 47
rect 132 46 133 52
rect 149 46 150 58
rect 152 46 153 58
rect 183 65 188 69
rect 179 59 180 65
rect 182 59 188 65
rect 189 49 190 54
rect 183 48 190 49
rect 192 48 194 54
rect 199 48 200 54
rect 202 48 203 54
rect 219 48 220 60
rect 222 48 223 60
rect 229 48 230 60
rect 232 48 233 60
<< ndcontact >>
rect 13 28 19 34
rect 53 25 59 34
rect 63 28 69 34
rect 83 28 89 34
rect 93 28 99 34
rect 103 28 109 34
rect 113 28 119 34
rect 143 25 149 34
rect 153 25 159 34
rect 173 24 178 28
rect 184 30 189 34
rect 194 32 199 36
rect 223 28 229 36
rect 183 13 188 17
<< pdcontact >>
rect 183 69 189 73
rect 13 46 19 52
rect 33 46 39 52
rect 53 46 59 58
rect 63 46 69 55
rect 83 46 89 52
rect 103 46 109 55
rect 113 46 119 52
rect 133 46 139 52
rect 143 46 149 58
rect 153 46 159 58
rect 173 59 179 65
rect 183 49 189 54
rect 194 48 199 54
rect 223 48 229 60
<< psubstratepcontact >>
rect 28 10 42 17
rect 91 10 105 17
rect 154 10 168 17
rect 194 10 208 17
rect 223 10 237 17
<< nsubstratencontact >>
rect 28 69 42 76
rect 91 69 105 76
rect 154 69 168 76
rect 194 69 208 76
rect 223 69 237 76
<< polysilicon >>
rect 10 19 12 67
rect 20 52 22 67
rect 30 52 32 67
rect 20 43 22 46
rect 30 43 32 46
rect 20 34 22 37
rect 30 34 32 37
rect 20 19 22 28
rect 30 19 32 28
rect 40 19 42 67
rect 50 55 52 67
rect 60 58 62 67
rect 70 63 72 67
rect 80 63 82 67
rect 50 43 52 46
rect 60 43 62 46
rect 70 43 72 46
rect 80 43 82 46
rect 50 34 52 37
rect 60 34 62 37
rect 70 34 72 37
rect 80 34 82 37
rect 50 19 52 28
rect 60 19 62 25
rect 70 19 72 20
rect 80 19 82 20
rect 90 19 92 67
rect 100 63 102 67
rect 100 55 102 58
rect 100 43 102 46
rect 100 34 102 37
rect 100 19 102 28
rect 110 19 112 67
rect 120 52 122 67
rect 130 52 132 67
rect 120 43 122 46
rect 130 43 132 46
rect 120 34 122 37
rect 130 34 132 37
rect 120 19 122 28
rect 130 19 132 28
rect 140 19 142 67
rect 150 58 152 67
rect 150 43 152 46
rect 150 34 152 37
rect 150 19 152 25
rect 160 19 162 67
rect 170 19 172 67
rect 180 65 182 68
rect 190 62 192 67
rect 200 63 202 67
rect 180 41 182 59
rect 190 54 192 57
rect 200 54 202 58
rect 190 45 192 48
rect 200 45 202 48
rect 180 25 182 37
rect 190 36 192 39
rect 200 36 202 39
rect 190 27 192 30
rect 200 26 202 32
rect 180 18 182 21
rect 190 19 192 22
rect 200 19 202 21
rect 210 19 212 67
rect 220 60 222 67
rect 230 60 232 67
rect 220 36 222 48
rect 230 45 232 48
rect 230 36 232 39
rect 220 25 222 28
rect 230 19 232 28
rect 240 19 242 67
<< polycontact >>
rect 18 37 24 43
rect 78 58 84 63
rect 48 37 53 43
rect 78 20 84 25
rect 98 58 104 63
rect 100 37 104 43
rect 118 37 124 43
rect 178 37 182 41
rect 228 39 234 45
rect 218 20 222 25
<< polypplus >>
rect 70 55 72 58
rect 80 55 82 58
<< polynplus >>
rect 20 28 22 30
rect 30 28 32 30
rect 70 25 72 28
rect 80 25 82 28
<< metal1 >>
rect 6 76 246 77
rect 6 69 28 76
rect 42 69 91 76
rect 105 69 154 76
rect 168 73 194 76
rect 168 69 183 73
rect 189 69 194 73
rect 208 69 223 76
rect 237 69 246 76
rect 13 52 19 69
rect 33 52 39 69
rect 53 58 59 69
rect 84 58 98 63
rect 113 55 119 69
rect 69 46 70 55
rect 13 37 18 43
rect 66 34 70 46
rect 83 34 89 40
rect 13 17 19 28
rect 69 28 70 34
rect 92 46 93 54
rect 109 52 119 55
rect 109 46 113 52
rect 133 52 139 69
rect 143 58 149 69
rect 168 59 173 65
rect 179 59 180 65
rect 159 46 164 58
rect 92 34 97 46
rect 157 45 164 46
rect 110 37 118 43
rect 157 39 159 45
rect 157 34 164 39
rect 92 28 93 34
rect 109 28 113 34
rect 92 25 99 28
rect 53 17 59 25
rect 84 20 99 25
rect 113 17 119 28
rect 159 25 164 34
rect 168 39 174 59
rect 223 60 229 69
rect 189 49 191 54
rect 173 34 174 39
rect 168 28 174 34
rect 189 30 191 34
rect 194 45 199 48
rect 194 39 228 45
rect 194 36 199 39
rect 143 17 149 25
rect 168 24 173 28
rect 225 17 229 28
rect 6 10 28 17
rect 42 10 91 17
rect 105 10 154 17
rect 168 13 183 17
rect 188 13 194 17
rect 168 10 194 13
rect 208 10 223 17
rect 237 10 246 17
rect 6 9 246 10
<< m2contact >>
rect 104 58 110 64
rect 7 37 13 43
rect 104 37 110 43
rect 213 20 218 25
<< pm12contact >>
rect 68 58 74 63
rect 28 37 34 43
rect 58 37 63 43
rect 128 37 134 43
rect 148 37 154 43
rect 68 20 74 25
rect 189 57 194 62
rect 198 58 203 63
rect 189 22 194 27
rect 198 21 203 26
<< pdm12contact >>
rect 23 47 29 53
rect 43 47 49 55
rect 73 46 79 52
rect 93 46 99 54
rect 123 47 129 53
rect 203 48 209 54
rect 213 48 219 60
rect 233 48 239 60
<< ndm12contact >>
rect 33 27 39 33
rect 43 27 49 33
rect 73 29 79 34
rect 133 27 139 33
rect 203 30 209 36
rect 213 29 219 36
rect 233 28 239 36
<< metal2 >>
rect 63 73 69 79
rect 7 43 13 71
rect 63 67 110 73
rect 104 64 110 67
rect 33 58 39 59
rect 7 26 13 37
rect 17 33 23 53
rect 74 58 99 62
rect 68 56 99 58
rect 33 43 39 52
rect 93 54 99 56
rect 49 47 58 53
rect 34 37 39 43
rect 52 33 58 47
rect 17 27 27 33
rect 49 27 58 33
rect 73 35 79 46
rect 104 43 110 58
rect 168 57 189 62
rect 168 39 173 57
rect 73 34 84 35
rect 79 29 84 34
rect 78 15 84 29
rect 104 26 110 37
rect 177 27 182 41
rect 203 45 209 48
rect 213 45 219 48
rect 203 39 219 45
rect 203 36 209 39
rect 213 36 219 39
rect 236 36 239 48
rect 177 22 189 27
rect 212 20 213 25
rect 212 15 218 20
rect 78 9 218 15
<< m3contact >>
rect 6 71 14 79
rect 33 52 39 58
rect 63 37 69 43
rect 27 27 33 33
rect 203 58 208 63
rect 117 47 123 53
rect 122 37 128 43
rect 143 37 148 43
rect 7 20 13 26
rect 62 20 68 26
rect 139 27 145 33
rect 223 36 236 48
rect 104 20 110 26
rect 203 21 208 26
<< m123contact >>
rect 43 37 48 43
rect 83 40 89 46
rect 159 39 164 45
rect 168 34 173 39
rect 177 41 182 46
rect 186 34 191 49
<< metal3 >>
rect 158 69 242 75
rect 123 47 145 53
rect 27 37 43 43
rect 69 40 83 43
rect 139 43 145 47
rect 158 45 164 69
rect 236 66 242 69
rect 89 40 122 43
rect 69 37 122 40
rect 139 37 143 43
rect 158 39 159 45
rect 177 58 203 63
rect 236 60 246 66
rect 177 46 182 58
rect 27 33 33 37
rect 139 33 145 37
rect 240 39 246 60
rect 168 26 173 34
rect 13 20 31 23
rect 68 20 104 26
rect 168 21 203 26
rect 7 17 31 20
rect 25 15 31 17
rect 6 7 14 13
rect 25 9 246 15
rect 237 7 246 9
<< m345contact >>
rect 32 58 39 65
<< metal5 >>
rect 6 58 32 65
rect 39 58 246 65
<< labels >>
rlabel nsubstratencontact 230 73 230 73 7 Vdd
rlabel metal5 7 62 7 62 3 y
rlabel m123contact 179 43 179 43 1 enable
rlabel metal1 194 13 194 13 1 Gnd
rlabel metal1 196 41 196 41 1 mux_out
rlabel metal2 206 43 206 43 1 D
rlabel m3contact 10 75 10 75 3 x
rlabel metal2 81 18 81 18 1 z
rlabel metal2 66 78 66 78 5 p
<< end >>
