magic
tech scmos
timestamp 1576137657
<< pwell >>
rect 6083 -8508 6125 -8485
rect 6083 -8527 6087 -8508
rect 6083 -8608 6125 -8527
<< metal1 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1543 13975 1569
rect -1773 1541 15766 1543
rect -1773 1529 15098 1541
rect -1773 1232 -1767 1529
rect -754 1232 15098 1529
rect -1773 1214 15098 1232
rect -1773 226 -1444 1214
rect 15425 1214 15766 1541
rect 15437 1197 15766 1214
rect -1773 -623 -1772 226
rect -1449 -623 -1444 226
rect -1773 -654 -1444 -623
rect -1216 657 14878 986
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -1336 -1441 -665
rect -3013 -1341 -1441 -1336
rect -1773 -15993 -1444 -1341
rect -1216 -15423 -887 657
rect 232 650 561 657
rect 14873 645 14878 657
rect 15437 868 15441 1197
rect 232 456 561 457
rect -667 127 14661 456
rect -666 -14873 -337 127
rect -116 -95 213 -94
rect 577 -95 14100 -94
rect -116 -423 14100 -95
rect -116 -14336 213 -423
rect 13771 -3679 14100 -423
rect 13756 -4525 14100 -3679
rect 10730 -5180 10840 -5153
rect 10870 -5153 10930 -5150
rect 10870 -5180 10952 -5153
rect 9731 -5532 9848 -5502
rect 10878 -5588 10905 -5180
rect 10730 -5618 10840 -5591
rect 10870 -5618 10930 -5588
rect 9701 -5934 9848 -5933
rect 9731 -5963 9848 -5934
rect 9731 -5964 9791 -5963
rect 10878 -6017 10905 -5618
rect 10730 -6047 10841 -6021
rect 10871 -6047 10931 -6017
rect 10730 -6048 10905 -6047
rect 9731 -6400 9848 -6370
rect 10878 -6452 10905 -6048
rect 10730 -6482 10835 -6455
rect 10865 -6482 10925 -6452
rect 9731 -6834 9848 -6804
rect 10878 -6886 10905 -6482
rect 10730 -6916 10828 -6889
rect 10858 -6916 10918 -6886
rect 6423 -7141 6448 -7117
rect 6490 -7141 7390 -7117
rect 6423 -7142 7390 -7141
rect 6514 -7174 6526 -7142
rect 6618 -7174 6630 -7142
rect 6722 -7174 6734 -7142
rect 6826 -7174 6838 -7142
rect 6930 -7174 6942 -7142
rect 7034 -7174 7046 -7142
rect 7138 -7176 7150 -7142
rect 7242 -7174 7254 -7142
rect 5306 -7429 5331 -7329
rect 5616 -7353 5783 -7341
rect 5795 -7353 5815 -7341
rect 5776 -7404 5788 -7353
rect 6426 -7404 6438 -7382
rect 5776 -7425 5789 -7404
rect 6426 -7425 6441 -7404
rect 5244 -7441 5268 -7429
rect 5280 -7441 5386 -7429
rect 5306 -7533 5331 -7441
rect 5776 -7445 5788 -7425
rect 6530 -7404 6542 -7382
rect 6634 -7404 6646 -7382
rect 6738 -7404 6750 -7382
rect 6842 -7404 6854 -7382
rect 6946 -7404 6958 -7382
rect 7050 -7404 7062 -7382
rect 7154 -7404 7166 -7382
rect 7285 -7404 7297 -7403
rect 7763 -7404 7784 -7156
rect 9731 -7268 9848 -7238
rect 10878 -7320 10905 -6916
rect 10730 -7350 10840 -7323
rect 10870 -7350 10930 -7320
rect 6483 -7425 7784 -7404
rect 5615 -7457 5775 -7445
rect 5787 -7457 5788 -7445
rect 5246 -7545 5270 -7533
rect 5282 -7545 5386 -7533
rect 5306 -7637 5331 -7545
rect 5776 -7549 5788 -7457
rect 5615 -7561 5766 -7549
rect 5778 -7561 5788 -7549
rect 5247 -7649 5271 -7637
rect 5283 -7649 5387 -7637
rect 5306 -7741 5331 -7649
rect 5776 -7653 5788 -7561
rect 8810 -7602 9068 -7594
rect 5616 -7665 5768 -7653
rect 5780 -7665 5788 -7653
rect 8810 -7662 8899 -7654
rect 5249 -7753 5273 -7741
rect 5285 -7753 5388 -7741
rect 5306 -7845 5331 -7753
rect 5776 -7757 5788 -7665
rect 8810 -7674 9067 -7666
rect 9075 -7674 9076 -7666
rect 9731 -7702 9848 -7672
rect 8810 -7734 8879 -7726
rect 8887 -7734 8927 -7726
rect 8810 -7746 9077 -7738
rect 10878 -7754 10905 -7350
rect 5616 -7769 5789 -7757
rect 5251 -7857 5275 -7845
rect 5287 -7857 5387 -7845
rect 5306 -7949 5331 -7857
rect 5776 -7861 5788 -7769
rect 10730 -7784 10834 -7757
rect 10864 -7784 10924 -7754
rect 8810 -7806 8879 -7798
rect 8810 -7818 9073 -7810
rect 5616 -7873 5788 -7861
rect 5249 -7961 5273 -7949
rect 5285 -7961 5386 -7949
rect 5306 -8053 5331 -7961
rect 5776 -7965 5788 -7873
rect 8810 -7878 8877 -7870
rect 8810 -7890 9075 -7882
rect 8810 -7950 8876 -7942
rect 8809 -7962 9077 -7954
rect 5616 -7977 5774 -7965
rect 5786 -7977 5788 -7965
rect 5245 -8065 5270 -8053
rect 5282 -8065 5392 -8053
rect 5306 -8157 5331 -8065
rect 5776 -8069 5788 -7977
rect 8810 -8022 8877 -8014
rect 8810 -8034 9076 -8026
rect 5616 -8081 5788 -8069
rect 8810 -8094 8885 -8086
rect 8810 -8106 9075 -8098
rect 9731 -8136 9848 -8106
rect 5258 -8169 5282 -8157
rect 5294 -8169 5386 -8157
rect 8810 -8166 8883 -8158
rect 10878 -8188 10905 -7784
rect 10730 -8218 10832 -8191
rect 10862 -8218 10922 -8188
rect 5783 -8346 5807 -8334
rect 5819 -8346 6766 -8334
rect 6027 -8378 6039 -8346
rect 6131 -8378 6143 -8346
rect 6235 -8378 6247 -8346
rect 6339 -8378 6351 -8346
rect 6443 -8378 6455 -8346
rect 6547 -8378 6559 -8346
rect 6651 -8378 6663 -8346
rect 6754 -8386 6766 -8346
rect 10100 -8429 10104 -8424
rect 9731 -8570 9848 -8540
rect 10878 -8570 10905 -8218
rect 5237 -8644 5261 -8632
rect 5273 -8633 6039 -8632
rect 6115 -8633 6127 -8608
rect 6219 -8633 6231 -8608
rect 6323 -8633 6335 -8608
rect 6427 -8633 6439 -8605
rect 6531 -8633 6543 -8608
rect 6635 -8633 6647 -8608
rect 6739 -8633 6751 -8608
rect 6844 -8633 6856 -8592
rect 5273 -8644 6856 -8633
rect 6027 -8645 6856 -8644
rect 6963 -9871 6990 -9743
rect 6963 -9925 6990 -9898
rect 7282 -10085 7309 -9743
rect 7398 -9884 7425 -9743
rect 7398 -9938 7425 -9911
rect 7282 -10139 7309 -10112
rect 7716 -10085 7743 -9743
rect 7831 -9886 7858 -9743
rect 7831 -9940 7858 -9913
rect 7716 -10139 7743 -10112
rect 8150 -10084 8177 -9743
rect 8264 -9888 8291 -9743
rect 8264 -9940 8291 -9915
rect 8584 -10089 8611 -9743
rect 8708 -9884 8735 -9743
rect 8708 -9938 8735 -9911
rect 9018 -10089 9045 -9743
rect 9150 -9884 9177 -9743
rect 9176 -9911 9177 -9884
rect 9150 -9938 9177 -9911
rect 8150 -10138 8177 -10111
rect 8610 -10116 8611 -10089
rect 9044 -10116 9045 -10089
rect 8584 -10142 8611 -10116
rect 9018 -10143 9045 -10116
rect 9452 -10089 9479 -9743
rect 9569 -9882 9596 -9743
rect 9569 -9936 9596 -9909
rect 9452 -10142 9479 -10116
rect 9886 -10089 9913 -9743
rect 10010 -9880 10037 -9743
rect 10036 -9907 10037 -9880
rect 10010 -9934 10037 -9907
rect 9886 -10143 9913 -10116
rect 10320 -10090 10347 -9743
rect 10320 -10144 10347 -10117
rect 13756 -14333 14085 -4525
rect -116 -14341 222 -14336
rect 582 -14341 13655 -14336
rect -116 -14658 13655 -14341
rect -116 -14665 222 -14658
rect 588 -14665 13655 -14658
rect 14323 -14871 14655 127
rect 14873 -1424 15202 645
rect 232 -14873 561 -14872
rect 866 -14873 14655 -14871
rect -666 -14876 14655 -14873
rect -666 -15202 14211 -14876
rect -664 -15211 14211 -15202
rect 14645 -15200 14655 -14876
rect 14870 -3055 15202 -1424
rect 14870 -14709 15199 -3055
rect 15437 -13974 15766 868
rect 15434 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 14870 -15053 14871 -14709
rect 15437 -14766 15766 -14654
rect 14645 -15211 14649 -15200
rect 14870 -15418 15199 -15053
rect 232 -15423 561 -15420
rect -1216 -15752 14778 -15423
rect 15521 -14799 15766 -14766
rect 15521 -15983 15646 -14799
rect 15437 -15989 15646 -15983
rect 10 -15993 661 -15992
rect 15437 -15993 15768 -15989
rect -1773 -15998 8414 -15993
rect -1773 -16081 14470 -15998
rect -1773 -16210 15766 -16081
rect -1773 -16315 14469 -16210
rect -1773 -16322 10 -16315
rect 661 -16322 14469 -16315
rect 7835 -16324 14469 -16322
rect 15753 -16324 15766 -16210
rect 7835 -16327 15766 -16324
rect 10 -17229 661 -16553
<< metal2 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1546 13975 1569
rect 240 1543 15763 1546
rect -1774 1541 15763 1543
rect -1774 1538 15098 1541
rect -1774 1529 13299 1538
rect -1774 1232 -1767 1529
rect -754 1232 13299 1529
rect -1774 1217 13299 1232
rect -1774 1214 890 1217
rect -1774 1211 -1445 1214
rect -1774 255 -1767 1211
rect -1456 255 -1445 1211
rect 13971 1217 15098 1538
rect 15425 1219 15436 1541
rect 15758 1219 15763 1541
rect 15425 1217 15763 1219
rect 15434 1197 15763 1217
rect -929 981 14512 982
rect -1774 226 -1445 255
rect -1774 -623 -1772 226
rect -1449 -623 -1445 226
rect -1774 -654 -1445 -623
rect -1217 814 14512 981
rect -1217 664 12407 814
rect 13092 664 14512 814
rect -1217 660 14512 664
rect 14852 660 14878 982
rect -1217 653 14878 660
rect -1217 652 896 653
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -670 -1441 -665
rect -1835 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -1835 -1336 -1441 -1331
rect -3013 -1341 -1441 -1336
rect -1774 -15992 -1445 -1341
rect -1217 -1544 -888 652
rect 15434 868 15441 1197
rect 14884 618 15213 645
rect -1217 -2224 -1047 -1544
rect -889 -2224 -888 -1544
rect -1217 -15428 -888 -2224
rect -667 444 876 457
rect -667 129 14649 444
rect -667 -14001 -339 129
rect 467 116 14649 129
rect 1720 -95 2049 -94
rect 2520 -95 14096 -93
rect -116 -422 14096 -95
rect -116 -423 3442 -422
rect -116 -424 222 -423
rect 582 -424 3442 -423
rect -116 -13100 213 -424
rect 13767 -1532 14096 -422
rect 13932 -2213 14096 -1532
rect 10729 -5417 10779 -5302
rect 10729 -5851 10768 -5736
rect 10729 -6285 10768 -6170
rect 10729 -6719 10768 -6604
rect 10729 -7154 10768 -7039
rect 10729 -7587 10768 -7472
rect 10729 -8021 10768 -7906
rect 10729 -8456 10768 -8341
rect -116 -13787 42 -13100
rect 200 -13787 213 -13100
rect -667 -14674 -482 -14001
rect -116 -14333 213 -13787
rect 13767 -13979 14096 -2213
rect 14095 -14312 14096 -13979
rect 13767 -14333 14096 -14312
rect 14321 -636 14649 116
rect 14321 -1321 14327 -636
rect 14499 -1321 14649 -636
rect -116 -14341 222 -14333
rect 582 -14341 13267 -14333
rect -116 -14347 13267 -14341
rect -116 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -116 -14662 13267 -14484
rect 13646 -14662 13655 -14333
rect 14321 -14517 14649 -1321
rect 14884 -13082 15213 272
rect 15028 -13769 15213 -13082
rect -667 -14883 -339 -14674
rect 14321 -14850 14327 -14517
rect 14884 -14709 15213 -13769
rect 14321 -14876 14649 -14850
rect -667 -15043 13336 -14883
rect 14002 -15043 14211 -14883
rect -667 -15211 14211 -15043
rect 14645 -15211 14649 -14876
rect 15212 -15053 15213 -14709
rect 14884 -15063 15213 -15053
rect 15212 -15398 15213 -15063
rect 14884 -15418 15213 -15398
rect -1217 -15609 14338 -15428
rect -1217 -15757 886 -15609
rect 1567 -15757 14338 -15609
rect 14772 -15757 14778 -15428
rect 15212 -15757 15213 -15418
rect 15434 -13972 15763 868
rect 15434 -14674 15436 -13972
rect 15747 -13974 15763 -13972
rect 15747 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 15747 -14674 15763 -14654
rect 15434 -14694 15763 -14674
rect 15434 -14766 15766 -14694
rect 15521 -14771 15766 -14766
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -14799 15766 -14771
rect 15644 -15986 15646 -14799
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16081 14470 -15993
rect 662 -16090 15766 -16081
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16210 15766 -16204
rect 662 -16313 14469 -16210
rect -1774 -16315 14469 -16313
rect -1774 -16321 10 -16315
rect -9 -16322 10 -16321
rect 661 -16321 14469 -16315
rect 15753 -16321 15766 -16210
rect 10 -17229 661 -16553
<< m123contact >>
rect 13308 1569 13962 1943
rect -1767 1232 -754 1529
rect 15098 1212 15425 1541
rect -1772 -623 -1449 226
rect -2255 -1336 -1835 -665
rect 14878 645 15219 991
rect 15441 868 15768 1197
rect 10840 -5180 10870 -5150
rect 9701 -5532 9731 -5502
rect 10840 -5618 10870 -5588
rect 9701 -5964 9731 -5934
rect 10841 -6047 10871 -6017
rect 9701 -6400 9731 -6370
rect 10835 -6482 10865 -6452
rect 9701 -6834 9731 -6804
rect 10828 -6916 10858 -6886
rect 6448 -7141 6490 -7117
rect 9701 -7268 9731 -7238
rect 5783 -7353 5795 -7341
rect 10840 -7350 10870 -7320
rect 6441 -7427 6483 -7403
rect 5268 -7441 5280 -7429
rect 5775 -7457 5787 -7445
rect 5270 -7545 5282 -7533
rect 5766 -7561 5778 -7549
rect 8488 -7602 8496 -7594
rect 9068 -7602 9076 -7594
rect 5271 -7649 5283 -7637
rect 5768 -7665 5780 -7653
rect 7642 -7660 7650 -7654
rect 8899 -7662 8907 -7654
rect 7402 -7672 7410 -7666
rect 8487 -7674 8495 -7668
rect 9067 -7674 9075 -7666
rect 9701 -7702 9731 -7672
rect 8879 -7734 8887 -7726
rect 5273 -7753 5285 -7741
rect 9077 -7746 9085 -7738
rect 10834 -7784 10864 -7754
rect 7591 -7804 7599 -7798
rect 8628 -7804 8636 -7798
rect 8879 -7806 8887 -7798
rect 9073 -7818 9081 -7810
rect 5275 -7857 5287 -7845
rect 8632 -7876 8640 -7870
rect 8877 -7878 8885 -7870
rect 8686 -7888 8694 -7882
rect 9075 -7890 9083 -7882
rect 8647 -7948 8655 -7942
rect 5273 -7961 5285 -7949
rect 8876 -7950 8884 -7942
rect 8683 -7960 8691 -7954
rect 9077 -7962 9085 -7954
rect 5774 -7977 5786 -7965
rect 8632 -8020 8640 -8014
rect 8877 -8022 8885 -8014
rect 9076 -8034 9084 -8026
rect 5270 -8065 5282 -8053
rect 8681 -8092 8689 -8086
rect 8885 -8094 8893 -8086
rect 8638 -8104 8646 -8098
rect 9075 -8106 9083 -8098
rect 9701 -8136 9731 -8106
rect 5282 -8169 5294 -8157
rect 8655 -8164 8663 -8158
rect 8883 -8166 8891 -8158
rect 10832 -8218 10862 -8188
rect 5807 -8346 5819 -8334
rect 9701 -8570 9731 -8540
rect 5261 -8644 5273 -8632
rect 6963 -9898 6990 -9871
rect 7398 -9911 7425 -9884
rect 7831 -9913 7858 -9886
rect 8264 -9915 8291 -9888
rect 8708 -9911 8735 -9884
rect 9149 -9911 9176 -9884
rect 9569 -9909 9596 -9882
rect 10009 -9907 10036 -9880
rect 7282 -10112 7309 -10085
rect 7716 -10112 7743 -10085
rect 8150 -10111 8177 -10084
rect 8583 -10116 8610 -10089
rect 9017 -10116 9044 -10089
rect 9452 -10116 9479 -10089
rect 9886 -10116 9913 -10089
rect 10320 -10117 10347 -10090
rect 13655 -14672 14099 -14333
rect 14211 -15222 14645 -14876
rect 14871 -15053 15212 -14709
rect 14778 -15764 15212 -15418
rect 15766 -14654 15975 -13974
rect 15434 -15983 15521 -14766
rect 15646 -15989 15768 -14799
rect 14470 -16081 15768 -15993
rect 10 -16553 661 -16315
rect 14469 -16324 15753 -16210
<< metal3 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1546 13975 1569
rect -1774 1541 15763 1546
rect -1774 1538 15098 1541
rect -1774 1529 13299 1538
rect -1774 1232 -1767 1529
rect -754 1232 13299 1529
rect -1774 1217 13299 1232
rect -1774 1211 -1445 1217
rect -1774 255 -1767 1211
rect -1456 255 -1445 1211
rect 13971 1217 15098 1538
rect 15425 1219 15436 1541
rect 15758 1219 15763 1541
rect 15425 1217 15763 1219
rect 15434 1197 15763 1217
rect -1774 226 -1445 255
rect -1774 -623 -1772 226
rect -1449 -623 -1445 226
rect -1774 -654 -1445 -623
rect -1224 982 1544 984
rect -1224 814 14512 982
rect -1224 664 12407 814
rect 13092 664 14512 814
rect -1224 660 14512 664
rect 14852 660 14878 982
rect -1224 655 14878 660
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -670 -1441 -665
rect -1835 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -1835 -1336 -1441 -1331
rect -3013 -1341 -1441 -1336
rect -1774 -15992 -1445 -1341
rect -1224 -1544 -895 655
rect 466 653 14878 655
rect 15434 868 15441 1197
rect 14884 618 15213 645
rect -667 444 1547 454
rect -667 125 14656 444
rect -1224 -2224 -1047 -1544
rect -1224 -15428 -895 -2224
rect -667 -14001 -338 125
rect 108 115 14656 125
rect -115 -101 2593 -94
rect -115 -423 14094 -101
rect -115 -13100 214 -423
rect 2416 -430 14094 -423
rect 13765 -1532 14094 -430
rect 13932 -2213 14094 -1532
rect 8399 -7628 8405 -7622
rect 8398 -7698 8405 -7694
rect -115 -13787 42 -13100
rect 200 -13787 214 -13100
rect -667 -14674 -482 -14001
rect -115 -14334 214 -13787
rect 13765 -13979 14094 -2213
rect 14327 -636 14656 115
rect 14499 -1321 14656 -636
rect 13765 -14333 14094 -14312
rect -115 -14347 13267 -14334
rect -115 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -115 -14663 13267 -14484
rect 13646 -14663 13655 -14334
rect 14327 -14517 14656 -1321
rect 14884 -13082 15213 272
rect 15028 -13769 15213 -13082
rect -667 -14889 -338 -14674
rect 14884 -14709 15213 -13769
rect 14327 -14876 14656 -14850
rect -667 -15043 13336 -14889
rect 14002 -15043 14211 -14889
rect -667 -15218 14211 -15043
rect 14645 -15218 14656 -14876
rect 15212 -15053 15213 -14709
rect 14884 -15063 15213 -15053
rect 15212 -15398 15213 -15063
rect 14884 -15418 15213 -15398
rect -1224 -15609 14338 -15428
rect -1224 -15757 886 -15609
rect 1567 -15757 14338 -15609
rect 14772 -15757 14778 -15428
rect 15212 -15757 15213 -15418
rect 15434 -13972 15763 868
rect 15434 -14674 15436 -13972
rect 15747 -13974 15763 -13972
rect 15747 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 15747 -14674 15763 -14654
rect 15434 -14694 15763 -14674
rect 15434 -14766 15766 -14694
rect 15521 -14771 15766 -14766
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -14799 15766 -14771
rect 15644 -15986 15646 -14799
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16081 14470 -15993
rect 662 -16090 15766 -16081
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16210 15766 -16204
rect 662 -16313 14469 -16210
rect -1774 -16315 14469 -16313
rect -1774 -16321 10 -16315
rect -9 -16322 10 -16321
rect 661 -16321 14469 -16315
rect 15753 -16321 15766 -16210
rect 10 -17229 661 -16553
<< m234contact >>
rect -1767 255 -1456 1211
rect 13299 1209 13971 1538
rect 15436 1219 15758 1541
rect 12407 664 13092 814
rect 14512 660 14852 987
rect -1816 -1331 -1462 -670
rect 14875 272 15216 618
rect -1047 -2224 -889 -1544
rect 13764 -2213 13932 -1532
rect 42 -13787 200 -13100
rect -482 -14674 -311 -14001
rect 14327 -1321 14499 -636
rect 13757 -14312 14095 -13979
rect 12441 -14484 13126 -14347
rect 13267 -14668 13646 -14333
rect 14872 -13769 15028 -13082
rect 14327 -14850 14665 -14517
rect 13336 -15043 14002 -14877
rect 14877 -15398 15212 -15063
rect 886 -15760 1567 -15609
rect 14338 -15757 14772 -15422
rect 15436 -14674 15747 -13972
rect 15529 -15986 15644 -14771
rect -7 -16313 662 -15992
rect 14468 -16204 15752 -16090
<< m4contact >>
rect 6466 -7156 6489 -7147
rect 6570 -7156 6593 -7147
rect 6674 -7156 6697 -7147
rect 6778 -7156 6801 -7147
rect 6882 -7156 6905 -7147
rect 6986 -7156 7009 -7147
rect 7090 -7156 7113 -7147
rect 7194 -7156 7217 -7147
rect 5373 -7401 5390 -7378
rect 6460 -7395 6484 -7380
rect 6564 -7395 6588 -7380
rect 6668 -7395 6692 -7380
rect 6772 -7395 6796 -7380
rect 6876 -7395 6900 -7380
rect 6980 -7395 7004 -7380
rect 7084 -7395 7108 -7380
rect 7188 -7395 7212 -7380
rect 5373 -7505 5390 -7482
rect 5373 -7609 5390 -7586
rect 8405 -7638 8412 -7622
rect 5373 -7713 5390 -7690
rect 5373 -7817 5390 -7794
rect 5373 -7921 5390 -7898
rect 5373 -8025 5390 -8002
rect 5373 -8129 5390 -8106
rect 6069 -8380 6093 -8356
rect 6173 -8380 6197 -8356
rect 6277 -8380 6301 -8356
rect 6381 -8380 6405 -8356
rect 6485 -8380 6509 -8356
rect 6589 -8380 6613 -8356
rect 6693 -8380 6717 -8356
rect 6797 -8380 6821 -8356
rect 6064 -8616 6087 -8604
rect 6168 -8616 6191 -8604
rect 6272 -8616 6295 -8604
rect 6376 -8616 6399 -8604
rect 6480 -8616 6503 -8604
rect 6584 -8616 6607 -8604
rect 6688 -8616 6711 -8604
rect 6792 -8616 6815 -8604
rect 7121 -8662 7143 -8645
rect 7555 -8662 7577 -8645
rect 7991 -8662 8013 -8645
rect 8424 -8662 8446 -8645
rect 8859 -8662 8881 -8645
rect 9294 -8662 9316 -8645
rect 9726 -8662 9748 -8645
rect 7050 -9791 7227 -9742
rect 7501 -9791 7678 -9742
rect 7921 -9791 8098 -9742
rect 8366 -9791 8543 -9742
rect 8802 -9791 8979 -9742
rect 9237 -9791 9414 -9742
rect 9662 -9791 9839 -9742
rect 10083 -9791 10260 -9742
<< metal4 >>
rect 13304 1549 13975 2669
rect 1879 1540 15436 1549
rect 15529 1541 15770 1549
rect 1879 1539 10833 1540
rect -1767 1537 10833 1539
rect -1767 1221 5718 1537
rect 5839 1224 10833 1537
rect 10954 1538 15436 1540
rect 10954 1224 13299 1538
rect 5839 1221 13299 1224
rect -1767 1220 13299 1221
rect -1767 1211 8012 1220
rect -1456 1210 8012 1211
rect -1456 255 -1438 1210
rect 13971 1220 15436 1538
rect 13971 1218 13975 1220
rect 15433 1219 15436 1220
rect 15758 1220 15770 1541
rect 15758 1219 15762 1220
rect -1767 -629 -1438 255
rect -1217 984 2672 989
rect -1217 976 14512 984
rect -1217 660 5184 976
rect 5305 975 14512 976
rect 5305 660 9714 975
rect -1767 -654 -1441 -629
rect -3013 -670 -1441 -654
rect -3013 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -3013 -1341 -1441 -1331
rect -1767 -1356 -1441 -1341
rect -1767 -10047 -1438 -1356
rect -1217 -1544 -888 660
rect 1910 659 9714 660
rect 9835 973 14512 975
rect 9835 823 12407 973
rect 13092 823 14512 973
rect 9835 814 14512 823
rect 9835 664 12407 814
rect 13092 664 14512 814
rect 9835 660 14512 664
rect 14852 660 15213 984
rect 9835 659 15213 660
rect 1910 655 15213 659
rect 14884 618 15213 655
rect -1217 -1546 -1047 -1544
rect -1217 -2226 -1215 -1546
rect -1057 -2224 -1047 -1546
rect -889 -2224 -888 -1544
rect -1057 -2226 -888 -2224
rect -1217 -9847 -888 -2226
rect -891 -9967 -888 -9847
rect -1443 -10167 -1438 -10047
rect -1767 -15992 -1438 -10167
rect -1217 -15415 -888 -9967
rect -667 451 2201 454
rect -667 444 14656 451
rect -667 443 9043 444
rect -667 127 7141 443
rect 7262 438 9043 443
rect 7262 127 8378 438
rect -667 125 8378 127
rect -667 -13991 -338 125
rect -322 122 8378 125
rect 8499 128 9043 438
rect 9164 128 14656 444
rect 8499 122 14656 128
rect -667 -14664 -663 -13991
rect -492 -14001 -338 -13991
rect -115 -94 6919 -87
rect -115 -102 14094 -94
rect -115 -103 8177 -102
rect -115 -416 6943 -103
rect -115 -13096 214 -416
rect 2735 -417 6943 -416
rect 7064 -417 8177 -103
rect 2735 -418 8177 -417
rect 8298 -104 14094 -102
rect 8298 -418 8842 -104
rect 2735 -420 8842 -418
rect 8963 -420 14094 -104
rect 2735 -423 14094 -420
rect 1188 -719 1527 -696
rect 846 -3560 869 -2769
rect 1504 -3225 1527 -719
rect 2092 -2755 2115 -695
rect 2972 -2524 2995 -723
rect 3866 -2182 3889 -724
rect 3866 -2205 4673 -2182
rect 2972 -2547 4419 -2524
rect 2092 -2778 4072 -2755
rect 1504 -3248 3569 -3225
rect 846 -3583 3011 -3560
rect 463 -3684 736 -3661
rect 713 -3948 736 -3684
rect 713 -3971 2547 -3948
rect 477 -4559 2137 -4536
rect 2114 -8106 2137 -4559
rect 2524 -8002 2547 -3971
rect 2988 -7898 3011 -3583
rect 3546 -7794 3569 -3248
rect 4049 -7690 4072 -2778
rect 4396 -7586 4419 -2547
rect 4650 -7482 4673 -2205
rect 4755 -7378 4778 -733
rect 5638 -2173 5670 -719
rect 5638 -2205 6396 -2173
rect 6364 -7147 6396 -2205
rect 6466 -7147 6485 -7146
rect 6570 -7147 6606 -709
rect 7391 -2151 7426 -708
rect 6674 -2186 7426 -2151
rect 6674 -7147 6709 -2186
rect 8263 -2548 8299 -680
rect 6778 -2584 8299 -2548
rect 6778 -7147 6814 -2584
rect 9186 -2901 9222 -658
rect 6883 -2937 9222 -2901
rect 6883 -7147 6919 -2937
rect 10076 -3226 10109 -655
rect 6987 -3259 10109 -3226
rect 6987 -7147 7020 -3259
rect 10948 -3471 10982 -663
rect 7091 -3505 10982 -3471
rect 7091 -7147 7125 -3505
rect 11831 -3793 11862 -637
rect 13765 -1530 14094 -423
rect 14327 -636 14656 122
rect 14499 -1321 14510 -636
rect 14327 -1323 14510 -1321
rect 13765 -1532 13945 -1530
rect 13932 -2213 13945 -1532
rect 7195 -3824 11862 -3793
rect 7195 -7147 7226 -3824
rect 6364 -7156 6466 -7147
rect 6364 -7165 6485 -7156
rect 6364 -7178 6466 -7165
rect 4755 -7401 5373 -7378
rect 6421 -7395 6460 -7387
rect 7270 -7383 8109 -7378
rect 7212 -7386 8109 -7383
rect 7212 -7391 7278 -7386
rect 4650 -7505 5373 -7482
rect 6421 -7550 6429 -7395
rect 6564 -7491 6572 -7395
rect 6673 -7448 6679 -7395
rect 6673 -7454 6707 -7448
rect 6701 -7477 6707 -7454
rect 6772 -7463 6780 -7395
rect 6876 -7450 6884 -7395
rect 6980 -7435 6988 -7395
rect 7085 -7418 7093 -7395
rect 7085 -7426 7869 -7418
rect 6980 -7443 7629 -7435
rect 6876 -7458 7389 -7450
rect 6772 -7471 7149 -7463
rect 6701 -7483 6907 -7477
rect 6564 -7499 6669 -7491
rect 6661 -7516 6669 -7499
rect 6901 -7518 6907 -7483
rect 7141 -7518 7149 -7471
rect 7381 -7528 7389 -7458
rect 7621 -7517 7629 -7443
rect 7861 -7518 7869 -7426
rect 8101 -7517 8109 -7386
rect 8412 -7562 8420 -7407
rect 8405 -7570 8420 -7562
rect 4396 -7609 5373 -7586
rect 8405 -7614 8413 -7570
rect 8405 -7622 8415 -7614
rect 4049 -7713 5373 -7690
rect 3546 -7817 5373 -7794
rect 5865 -7849 5869 -7841
rect 2988 -7921 5373 -7898
rect 2524 -8025 5373 -8002
rect 2114 -8129 5373 -8106
rect 5980 -8347 5989 -8238
rect 5980 -8356 6093 -8347
rect 6183 -8356 6190 -8241
rect 6354 -8260 6363 -8241
rect 6287 -8269 6363 -8260
rect 6287 -8356 6296 -8269
rect 6416 -8334 6423 -8241
rect 6660 -8292 6669 -8241
rect 6390 -8341 6423 -8334
rect 6496 -8301 6669 -8292
rect 6390 -8356 6397 -8341
rect 6496 -8356 6505 -8301
rect 6720 -8318 6729 -8237
rect 6600 -8327 6729 -8318
rect 6600 -8356 6609 -8327
rect 6901 -8333 6909 -8236
rect 6705 -8341 6909 -8333
rect 6705 -8356 6713 -8341
rect 6961 -8357 6969 -8236
rect 8314 -8263 8323 -7704
rect 6821 -8365 6969 -8357
rect 7124 -8272 8323 -8263
rect 6167 -8616 6168 -8615
rect 6191 -8616 6192 -8615
rect 6063 -12122 6088 -8616
rect -115 -13778 -111 -13096
rect 28 -13100 214 -13096
rect 28 -13778 42 -13100
rect -115 -13787 42 -13778
rect 200 -13787 214 -13100
rect -492 -14664 -482 -14001
rect -667 -14674 -482 -14664
rect -115 -14334 214 -13787
rect 2116 -12147 6088 -12122
rect 2116 -14244 2141 -12147
rect 6167 -12316 6192 -8616
rect 2975 -12341 6192 -12316
rect 6271 -8616 6272 -8614
rect 6295 -8616 6296 -8614
rect 2975 -14244 3000 -12341
rect 6271 -12458 6296 -8616
rect 3820 -12483 6296 -12458
rect 6399 -8616 6401 -8612
rect 3820 -14221 3845 -12483
rect 6376 -12629 6401 -8616
rect 4789 -12654 6401 -12629
rect 6479 -8616 6480 -8613
rect 6503 -8616 6504 -8613
rect 4789 -14217 4814 -12654
rect 6479 -12830 6504 -8616
rect 5650 -12855 6504 -12830
rect 6583 -8616 6584 -8613
rect 6607 -8616 6608 -8613
rect 5650 -14192 5675 -12855
rect 6583 -14194 6608 -8616
rect 6687 -8616 6688 -8613
rect 6711 -8616 6712 -8613
rect 6687 -13481 6712 -8616
rect 6791 -8616 6792 -8615
rect 6815 -8616 6816 -8615
rect 6791 -13286 6816 -8616
rect 7124 -8645 7133 -8272
rect 8314 -8273 8323 -8272
rect 8745 -7778 8749 -7769
rect 8327 -8291 8336 -7783
rect 7566 -8300 8336 -8291
rect 8747 -7850 8749 -7841
rect 7566 -8645 7575 -8300
rect 8340 -8337 8349 -7852
rect 8396 -7922 8410 -7914
rect 8402 -7942 8410 -7922
rect 8747 -7926 8749 -7917
rect 8002 -8346 8349 -8337
rect 8353 -8337 8362 -7954
rect 8366 -7995 8399 -7986
rect 8746 -7994 8749 -7985
rect 8366 -8318 8375 -7995
rect 8379 -8066 8400 -8057
rect 8379 -8292 8388 -8066
rect 8392 -8275 8401 -8139
rect 8392 -8284 9065 -8275
rect 8379 -8301 8954 -8292
rect 8366 -8327 8872 -8318
rect 8353 -8346 8435 -8337
rect 8002 -8645 8011 -8346
rect 8426 -8645 8435 -8346
rect 8863 -8645 8872 -8327
rect 8945 -8578 8954 -8301
rect 9056 -8506 9065 -8284
rect 9056 -8515 9557 -8506
rect 8945 -8587 9302 -8578
rect 9293 -8645 9302 -8587
rect 9293 -8657 9294 -8645
rect 9548 -8657 9557 -8515
rect 9548 -8662 9726 -8657
rect 9548 -8666 9734 -8662
rect 13521 -9791 13563 -9744
rect 7110 -9835 7156 -9791
rect 7563 -9832 7609 -9791
rect 7112 -12792 7156 -9835
rect 7564 -12452 7605 -9832
rect 7986 -9833 8032 -9791
rect 8431 -9832 8477 -9791
rect 8876 -9832 8922 -9791
rect 7986 -12168 8028 -9833
rect 8436 -11880 8477 -9832
rect 8881 -11575 8922 -9832
rect 9318 -9832 9364 -9791
rect 9761 -9832 9807 -9791
rect 9318 -11108 9359 -9832
rect 9766 -10717 9807 -9832
rect 10166 -9833 13563 -9791
rect 9766 -10758 13535 -10717
rect 9318 -11149 13491 -11108
rect 8881 -11616 13041 -11575
rect 8436 -11921 11864 -11880
rect 7986 -12210 11098 -12168
rect 7986 -12221 8028 -12210
rect 7564 -12493 10229 -12452
rect 7112 -12836 9200 -12792
rect 6791 -13311 8340 -13286
rect 6687 -13506 7470 -13481
rect 7445 -14196 7470 -13506
rect 8315 -14190 8340 -13311
rect 9156 -14159 9200 -12836
rect 10188 -14135 10229 -12493
rect 11056 -14152 11098 -12210
rect 11823 -14147 11864 -11921
rect 13000 -12501 13041 -11616
rect 13450 -11629 13491 -11149
rect 13450 -11670 13531 -11629
rect 13000 -12542 13544 -12501
rect 13765 -13979 14094 -2213
rect -115 -14346 13267 -14334
rect -115 -14662 6943 -14346
rect 7064 -14347 13267 -14346
rect 7064 -14348 12441 -14347
rect 7064 -14662 8178 -14348
rect -115 -14663 8178 -14662
rect 8299 -14663 8842 -14348
rect 8963 -14484 12441 -14348
rect 13126 -14484 13267 -14347
rect 8963 -14532 13267 -14484
rect 8963 -14663 12447 -14532
rect 13132 -14663 13267 -14532
rect 13765 -14334 14094 -14312
rect 13646 -14663 14094 -14334
rect 14327 -14517 14656 -1323
rect 14884 -9854 15213 272
rect 15207 -9971 15213 -9854
rect 14884 -13082 15213 -9971
rect 15028 -13761 15035 -13082
rect 15212 -13761 15213 -13082
rect 15028 -13769 15213 -13761
rect -667 -14882 -338 -14674
rect -667 -14899 13336 -14882
rect -667 -15211 7138 -14899
rect 7259 -15211 8375 -14899
rect 8496 -14900 13336 -14899
rect 8496 -15211 9041 -14900
rect 9162 -15043 13336 -14900
rect 14327 -14882 14656 -14850
rect 14002 -15043 14656 -14882
rect 9162 -15064 14656 -15043
rect 14884 -15063 15213 -13769
rect 9162 -15211 13341 -15064
rect 14007 -15211 14656 -15064
rect 15212 -15398 15213 -15063
rect 14884 -15415 15213 -15398
rect -1217 -15421 15213 -15415
rect -1217 -15598 886 -15421
rect 1567 -15422 15213 -15421
rect 1567 -15425 14338 -15422
rect 1567 -15437 10834 -15425
rect 1567 -15438 9716 -15437
rect 1567 -15598 5183 -15438
rect -1217 -15609 5183 -15598
rect -1217 -15744 886 -15609
rect 1567 -15744 5183 -15609
rect 5304 -15744 9716 -15438
rect 9837 -15741 10834 -15437
rect 10955 -15741 14338 -15425
rect 9837 -15744 14338 -15741
rect 14772 -15744 15213 -15422
rect 15433 -10053 15762 1219
rect 15433 -10170 15436 -10053
rect 15433 -13972 15762 -10170
rect 15433 -14674 15436 -13972
rect 15747 -13974 15762 -13972
rect 15747 -14654 16673 -13974
rect 15747 -14674 15762 -14654
rect 15433 -14694 15762 -14674
rect 15433 -14771 15766 -14694
rect 15433 -15986 15529 -14771
rect 15644 -15986 15766 -14771
rect 15433 -15989 15766 -15986
rect 15433 -15992 15768 -15989
rect -1788 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16005 15766 -15993
rect 662 -16313 5718 -16005
rect -1788 -16321 5718 -16313
rect 5839 -16007 15766 -16005
rect 5839 -16321 10836 -16007
rect -9 -16322 661 -16321
rect 10 -17229 661 -16322
rect 10957 -16016 15766 -16007
rect 10957 -16063 11215 -16016
rect 11336 -16063 15766 -16016
rect 10957 -16090 15766 -16063
rect 10957 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 10957 -16321 15766 -16204
<< m345contact >>
rect 6490 -7141 6532 -7117
rect 10870 -5180 10900 -5150
rect 9626 -5342 9649 -5318
rect 10729 -5417 10779 -5302
rect 9731 -5532 9761 -5502
rect 10870 -5618 10900 -5588
rect 9626 -5776 9649 -5752
rect 10729 -5851 10768 -5736
rect 9731 -5964 9761 -5934
rect 10871 -6047 10901 -6017
rect 9626 -6210 9649 -6186
rect 7563 -6284 7660 -6254
rect 10729 -6285 10768 -6170
rect 9731 -6400 9761 -6370
rect 10865 -6482 10895 -6452
rect 9626 -6644 9649 -6620
rect 10729 -6719 10768 -6604
rect 9731 -6834 9761 -6804
rect 10858 -6916 10888 -6886
rect 9626 -7078 9649 -7054
rect 10729 -7154 10768 -7039
rect 9731 -7268 9761 -7238
rect 5771 -7353 5783 -7341
rect 10870 -7350 10900 -7320
rect 7578 -7373 7600 -7364
rect 5614 -7407 5642 -7383
rect 5256 -7441 5268 -7429
rect 5763 -7457 5775 -7445
rect 5614 -7511 5642 -7487
rect 5258 -7545 5270 -7533
rect 5754 -7561 5766 -7549
rect 6483 -7428 6525 -7404
rect 9626 -7512 9649 -7488
rect 5614 -7615 5642 -7591
rect 10729 -7587 10768 -7472
rect 8496 -7602 8504 -7594
rect 9060 -7602 9068 -7594
rect 5259 -7649 5271 -7637
rect 5756 -7665 5768 -7653
rect 7650 -7660 7658 -7654
rect 8891 -7662 8899 -7654
rect 7410 -7672 7418 -7666
rect 8495 -7674 8503 -7668
rect 9059 -7674 9067 -7666
rect 5614 -7719 5642 -7695
rect 5261 -7753 5273 -7741
rect 5614 -7823 5642 -7799
rect 7599 -7804 7607 -7798
rect 5263 -7857 5275 -7845
rect 5614 -7927 5642 -7903
rect 5261 -7961 5273 -7949
rect 5762 -7977 5774 -7965
rect 5614 -8031 5642 -8007
rect 5258 -8065 5270 -8053
rect 5614 -8135 5642 -8111
rect 5270 -8169 5282 -8157
rect 5795 -8346 5807 -8334
rect 8405 -7710 8412 -7694
rect 9731 -7702 9761 -7672
rect 8871 -7734 8879 -7726
rect 9069 -7746 9077 -7738
rect 5249 -8644 5261 -8632
rect 8405 -7783 8412 -7768
rect 10864 -7784 10894 -7754
rect 8636 -7804 8644 -7798
rect 8871 -7806 8879 -7798
rect 9065 -7818 9073 -7810
rect 8640 -7876 8648 -7870
rect 8869 -7878 8877 -7870
rect 8694 -7888 8702 -7882
rect 9067 -7890 9075 -7882
rect 8655 -7948 8663 -7942
rect 8868 -7950 8876 -7942
rect 9626 -7946 9649 -7922
rect 8691 -7960 8699 -7954
rect 9069 -7962 9077 -7954
rect 8640 -8020 8648 -8014
rect 8869 -8022 8877 -8014
rect 10729 -8021 10768 -7906
rect 9068 -8034 9076 -8026
rect 8689 -8092 8697 -8086
rect 8877 -8094 8885 -8086
rect 8646 -8104 8654 -8098
rect 9067 -8106 9075 -8098
rect 9731 -8136 9761 -8106
rect 8663 -8164 8671 -8158
rect 8875 -8166 8883 -8158
rect 10862 -8218 10892 -8188
rect 9626 -8380 9649 -8356
rect 10729 -8456 10768 -8341
rect 9731 -8570 9761 -8540
rect 6963 -9925 6990 -9898
rect 7398 -9938 7425 -9911
rect 7282 -10139 7309 -10112
rect 7831 -9940 7858 -9913
rect 7716 -10139 7743 -10112
rect 8264 -9942 8291 -9915
rect 8150 -10138 8177 -10111
rect 8708 -9938 8735 -9911
rect 8583 -10143 8610 -10116
rect 9149 -9938 9176 -9911
rect 9017 -10143 9044 -10116
rect 9569 -9936 9596 -9909
rect 9452 -10143 9479 -10116
rect 10009 -9934 10036 -9907
rect 9886 -10143 9913 -10116
rect 10320 -10144 10347 -10117
<< m5contact >>
rect -1219 -9967 -891 -9847
rect -1771 -10167 -1443 -10047
rect 2092 -695 2115 -672
rect 1165 -719 1188 -696
rect 846 -2769 869 -2746
rect 2972 -723 2995 -700
rect 3866 -724 3889 -701
rect 4755 -733 4778 -710
rect 440 -3684 463 -3661
rect 454 -4559 477 -4536
rect 5638 -719 5670 -687
rect 6570 -709 6606 -673
rect 7391 -708 7426 -673
rect 8263 -680 8299 -644
rect 9186 -658 9222 -622
rect 10076 -655 10109 -622
rect 10948 -663 10982 -629
rect 11831 -637 11862 -606
rect 8412 -7407 8420 -7399
rect 8749 -7638 8758 -7625
rect 8314 -7704 8323 -7695
rect 5847 -7851 5865 -7839
rect 8749 -7710 8758 -7697
rect 2116 -14269 2141 -14244
rect 2975 -14269 3000 -14244
rect 3820 -14246 3845 -14221
rect 5650 -14217 5675 -14192
rect 8327 -7783 8336 -7770
rect 8749 -7782 8758 -7769
rect 8340 -7852 8349 -7843
rect 8401 -7852 8410 -7843
rect 8749 -7854 8758 -7841
rect 8749 -7926 8758 -7913
rect 8353 -7954 8362 -7945
rect 8402 -7950 8410 -7942
rect 8749 -7998 8758 -7985
rect 8749 -8070 8758 -8057
rect 8749 -8142 8758 -8129
rect 13521 -9744 13563 -9702
rect 13535 -10758 13576 -10717
rect 4789 -14242 4814 -14217
rect 6583 -14219 6608 -14194
rect 7445 -14221 7470 -14196
rect 8315 -14215 8340 -14190
rect 9156 -14203 9200 -14159
rect 10188 -14176 10229 -14135
rect 11056 -14194 11098 -14152
rect 13531 -11670 13572 -11629
rect 13544 -12542 13585 -12501
rect 11823 -14188 11864 -14147
rect 14877 -9971 15207 -9854
rect 15436 -10170 15766 -10053
<< metal5 >>
rect 1165 -696 1188 2050
rect 2092 -672 2115 2064
rect 2972 -700 2995 2064
rect 3866 -701 3889 2054
rect 4755 -710 4778 2054
rect 5639 -687 5670 2010
rect 6573 -673 6604 2014
rect 7394 -673 7425 2031
rect 8098 -613 8129 2071
rect 9364 -591 9395 2022
rect 8098 -644 8295 -613
rect 9186 -622 9395 -591
rect 10076 -622 10107 2039
rect 11090 -598 11121 2116
rect 10948 -629 11121 -598
rect 11831 -606 11862 2080
rect 12407 973 13089 2672
rect 12407 661 13089 823
rect 14325 -1320 14510 -640
rect 14657 -1320 16677 -640
rect -3000 -2224 -1215 -1549
rect -1057 -2224 -893 -1549
rect 13759 -2210 13945 -1533
rect 14102 -2210 16674 -1533
rect -2392 -2769 846 -2745
rect 13311 -2811 16033 -2766
rect -2443 -3684 440 -3660
rect -2411 -4559 454 -4536
rect -2411 -4560 465 -4559
rect 9446 -5341 9626 -5328
rect -2372 -5451 7598 -5429
rect 7576 -6254 7598 -5451
rect 9446 -5998 9459 -5341
rect 13311 -5339 13356 -2811
rect 10779 -5384 13356 -5339
rect 13497 -3706 16043 -3661
rect 9123 -6011 9459 -5998
rect 9483 -5776 9626 -5766
rect 9483 -5779 9634 -5776
rect 5812 -7054 6289 -7001
rect 5812 -7089 7130 -7054
rect 6201 -7117 7130 -7089
rect 6201 -7141 6490 -7117
rect 6532 -7141 7130 -7117
rect 6201 -7142 7130 -7141
rect 5186 -7242 5213 -7154
rect 5301 -7242 6089 -7154
rect 6001 -7404 6089 -7242
rect 7581 -7398 7594 -7373
rect 7581 -7399 8420 -7398
rect 5627 -7462 5635 -7407
rect 6001 -7428 6483 -7404
rect 6525 -7428 7142 -7404
rect 7581 -7407 8412 -7399
rect 7581 -7411 8420 -7407
rect 5627 -7470 5720 -7462
rect 5630 -7567 5641 -7511
rect 5630 -7578 5694 -7567
rect 5632 -7630 5640 -7615
rect 5632 -7638 5657 -7630
rect 5627 -7783 5635 -7719
rect 5649 -7757 5657 -7638
rect 5683 -7727 5694 -7578
rect 5712 -7684 5720 -7470
rect 6001 -7492 7142 -7428
rect 9123 -7625 9136 -6011
rect 9483 -6321 9496 -5779
rect 13497 -5763 13542 -3706
rect 10768 -5808 13542 -5763
rect 13613 -4590 16047 -4545
rect 8758 -7638 9136 -7625
rect 9162 -6334 9496 -6321
rect 9540 -6210 9626 -6198
rect 9540 -6211 9637 -6210
rect 5712 -7692 5812 -7684
rect 5683 -7738 5775 -7727
rect 5649 -7765 5747 -7757
rect 5627 -7791 5723 -7783
rect 5623 -7889 5631 -7823
rect 5623 -7897 5696 -7889
rect 5642 -7923 5670 -7918
rect 5632 -8064 5640 -8031
rect 5665 -8051 5670 -7923
rect 5688 -7942 5696 -7897
rect 5715 -7905 5723 -7791
rect 5739 -7870 5747 -7765
rect 5764 -7841 5775 -7738
rect 5804 -7769 5812 -7692
rect 8323 -7704 8405 -7695
rect 9162 -7697 9175 -6334
rect 9540 -6647 9553 -6211
rect 13613 -6213 13658 -4590
rect 10768 -6258 13658 -6213
rect 14141 -5456 16052 -5411
rect 8758 -7710 9175 -7697
rect 9192 -6660 9553 -6647
rect 9619 -6644 9626 -6622
rect 5804 -7777 5866 -7769
rect 8336 -7783 8405 -7770
rect 9192 -7769 9205 -6660
rect 9619 -6960 9632 -6644
rect 14141 -6623 14186 -5456
rect 10768 -6668 14186 -6623
rect 14710 -6362 16030 -6317
rect 8758 -7782 9205 -7769
rect 9244 -6973 9632 -6960
rect 5764 -7851 5847 -7841
rect 9244 -7841 9257 -6973
rect 9620 -7078 9626 -7055
rect 9620 -7281 9633 -7078
rect 14710 -7071 14755 -6362
rect 10768 -7116 14755 -7071
rect 15270 -7223 16087 -7178
rect 5865 -7849 5872 -7841
rect 5764 -7852 5849 -7851
rect 8349 -7852 8401 -7843
rect 8758 -7854 9257 -7841
rect 9288 -7294 9633 -7281
rect 5739 -7878 5866 -7870
rect 5715 -7913 5866 -7905
rect 9288 -7913 9301 -7294
rect 9618 -7512 9626 -7489
rect 9618 -7602 9631 -7512
rect 15270 -7519 15315 -7223
rect 10768 -7564 15315 -7519
rect 8758 -7914 8785 -7913
rect 8817 -7914 9301 -7913
rect 8758 -7926 9301 -7914
rect 9322 -7615 9631 -7602
rect 5688 -7950 5866 -7942
rect 8362 -7950 8402 -7942
rect 8362 -7954 8371 -7950
rect 9322 -7985 9335 -7615
rect 9622 -7946 9626 -7932
rect 9622 -7952 9635 -7946
rect 8825 -7988 9335 -7985
rect 8758 -7998 9335 -7988
rect 9363 -7965 9635 -7952
rect 5665 -8056 5865 -8051
rect 9363 -8057 9376 -7965
rect 10768 -8005 16061 -7960
rect 5632 -8072 5865 -8064
rect 8820 -8069 9376 -8057
rect 8758 -8070 9376 -8069
rect 8749 -8082 8833 -8070
rect 5666 -8113 5866 -8100
rect 5642 -8126 5679 -8113
rect 8811 -8141 9376 -8129
rect 8758 -8142 9376 -8141
rect 8749 -8154 8824 -8142
rect 8646 -8156 8653 -8154
rect 9363 -8350 9376 -8142
rect 9363 -8356 9641 -8350
rect 9363 -8363 9626 -8356
rect 10768 -8422 15323 -8377
rect 15278 -8972 15323 -8422
rect 15278 -9017 16047 -8972
rect 13563 -9744 16043 -9703
rect -891 -9854 15204 -9848
rect -891 -9898 14877 -9854
rect -891 -9925 6963 -9898
rect 6990 -9907 14877 -9898
rect 6990 -9909 10009 -9907
rect 6990 -9911 9569 -9909
rect 6990 -9925 7398 -9911
rect -891 -9938 7398 -9925
rect 7425 -9913 8708 -9911
rect 7425 -9938 7831 -9913
rect -891 -9940 7831 -9938
rect 7858 -9915 8708 -9913
rect 7858 -9940 8264 -9915
rect -891 -9942 8264 -9940
rect 8291 -9938 8708 -9915
rect 8735 -9938 9149 -9911
rect 9176 -9936 9569 -9911
rect 9596 -9934 10009 -9909
rect 10036 -9934 14877 -9907
rect 9596 -9936 14877 -9934
rect 9176 -9938 14877 -9936
rect 8291 -9942 14877 -9938
rect -891 -9967 14877 -9942
rect -1217 -9968 14877 -9967
rect -1775 -10167 -1771 -10049
rect -1443 -10053 15766 -10049
rect -1443 -10111 15436 -10053
rect -1443 -10112 8150 -10111
rect -1443 -10139 7282 -10112
rect 7309 -10139 7716 -10112
rect 7743 -10138 8150 -10112
rect 8177 -10116 15436 -10111
rect 8177 -10138 8583 -10116
rect 7743 -10139 8583 -10138
rect -1443 -10143 8583 -10139
rect 8610 -10143 9017 -10116
rect 9044 -10143 9452 -10116
rect 9479 -10143 9886 -10116
rect 9913 -10117 15436 -10116
rect 9913 -10143 10320 -10117
rect -1443 -10144 10320 -10143
rect 10347 -10144 15436 -10117
rect -1443 -10167 15436 -10144
rect -1775 -10169 15436 -10167
rect 13576 -10758 16057 -10717
rect 13571 -11629 16043 -11628
rect 13572 -11669 16043 -11629
rect 13585 -12542 16028 -12501
rect -3003 -13778 -111 -13096
rect 28 -13778 209 -13096
rect 14870 -13761 15035 -13086
rect 15212 -13761 16670 -13086
rect 14870 -13764 16670 -13761
rect -3003 -13787 209 -13778
rect -3009 -14664 -663 -13998
rect -492 -14664 -323 -13998
rect -3009 -14672 -323 -14664
rect 886 -15421 1565 -15415
rect 886 -17232 1565 -15598
rect 2116 -16694 2141 -14269
rect 2975 -16632 3000 -14269
rect 3820 -16730 3845 -14246
rect 4789 -16678 4814 -14242
rect 5650 -16683 5675 -14217
rect 6583 -16673 6608 -14219
rect 7445 -16642 7470 -14221
rect 8315 -16639 8340 -14215
rect 9158 -14806 9199 -14203
rect 9157 -14847 9340 -14806
rect 9158 -15217 9162 -15216
rect 9299 -15270 9340 -14847
rect 9158 -15311 9340 -15270
rect 9158 -16714 9199 -15311
rect 10188 -16632 10229 -14176
rect 11057 -14231 11098 -14194
rect 11061 -16666 11098 -14231
rect 11823 -16656 11864 -14188
rect 12444 -14532 13130 -14343
rect 12444 -14669 12447 -14532
rect 12444 -17227 13130 -14669
rect 13339 -15064 14003 -14871
rect 13339 -15230 13341 -15064
rect 13339 -17237 14003 -15230
<< m456contact >>
rect 5184 660 5305 976
rect 5718 1221 5839 1537
rect 7141 127 7262 443
rect 6943 -417 7064 -103
rect 8378 122 8499 438
rect 9043 128 9164 444
rect 8177 -418 8298 -102
rect 8842 -420 8963 -104
rect 9714 659 9835 975
rect 10833 1224 10954 1540
rect 12407 823 13092 973
rect 14510 -1323 14657 -636
rect -1215 -2226 -1057 -1546
rect 13945 -2213 14102 -1530
rect -111 -13778 28 -13096
rect 15035 -13761 15212 -13082
rect -663 -14664 -492 -13991
rect 886 -15598 1567 -15421
rect 5183 -15754 5304 -15438
rect 5718 -16321 5839 -16005
rect 6943 -14662 7064 -14346
rect 7138 -15215 7259 -14899
rect 8178 -14664 8299 -14348
rect 8842 -14664 8963 -14348
rect 8375 -15215 8496 -14899
rect 9041 -15216 9162 -14900
rect 9716 -15753 9837 -15437
rect 10836 -16323 10957 -16007
rect 12447 -14669 13132 -14532
rect 13341 -15230 14007 -15064
<< m6contact >>
rect 10900 -5180 10930 -5150
rect 9761 -5532 9791 -5502
rect 10900 -5618 10930 -5588
rect 5724 -7089 5812 -7001
rect 5213 -7242 5301 -7154
rect 5759 -7353 5771 -7341
rect 5244 -7441 5256 -7429
rect 5751 -7457 5763 -7445
rect 5246 -7545 5258 -7533
rect 5247 -7649 5259 -7637
rect 5249 -7753 5261 -7741
rect 5742 -7561 5754 -7549
rect 8504 -7602 8512 -7594
rect 9052 -7602 9060 -7594
rect 9761 -5964 9791 -5934
rect 10901 -6047 10931 -6017
rect 5744 -7665 5756 -7653
rect 7658 -7662 7666 -7654
rect 8883 -7662 8891 -7654
rect 7418 -7674 7426 -7666
rect 8503 -7676 8511 -7668
rect 9051 -7674 9059 -7666
rect 5251 -7857 5263 -7845
rect 5249 -7961 5261 -7949
rect 5246 -8065 5258 -8053
rect 9761 -6400 9791 -6370
rect 10895 -6482 10925 -6452
rect 8863 -7734 8871 -7726
rect 9061 -7746 9069 -7738
rect 9761 -6834 9791 -6804
rect 10888 -6916 10918 -6886
rect 7607 -7806 7615 -7798
rect 8644 -7806 8652 -7798
rect 8863 -7806 8871 -7798
rect 9057 -7818 9065 -7810
rect 9761 -7268 9791 -7238
rect 8648 -7878 8656 -7870
rect 8861 -7878 8869 -7870
rect 8702 -7890 8710 -7882
rect 9059 -7890 9067 -7882
rect 10900 -7350 10930 -7320
rect 8663 -7950 8671 -7942
rect 8860 -7950 8868 -7942
rect 8699 -7962 8707 -7954
rect 9061 -7962 9069 -7954
rect 5750 -7977 5762 -7965
rect 9761 -7702 9791 -7672
rect 10894 -7784 10924 -7754
rect 8648 -8022 8656 -8014
rect 8861 -8022 8869 -8014
rect 9060 -8034 9068 -8026
rect 8697 -8094 8705 -8086
rect 8869 -8094 8877 -8086
rect 8654 -8106 8662 -8098
rect 9059 -8106 9067 -8098
rect 9761 -8136 9791 -8106
rect 5258 -8169 5270 -8157
rect 8671 -8166 8679 -8158
rect 8867 -8166 8875 -8158
rect 5783 -8346 5795 -8334
rect 10892 -8218 10922 -8188
rect 9761 -8570 9791 -8540
rect 5237 -8644 5249 -8632
<< metal6 >>
rect 10836 1540 10956 1541
rect 5839 1221 5841 1517
rect 10954 1224 10956 1540
rect 5305 660 5307 948
rect -3000 -2224 -1215 -1549
rect -1057 -2224 -893 -1549
rect 5187 -7154 5307 660
rect 5187 -7242 5213 -7154
rect 5301 -7242 5307 -7154
rect 5187 -7429 5307 -7242
rect 5187 -7441 5244 -7429
rect 5256 -7441 5307 -7429
rect 5187 -7533 5307 -7441
rect 5187 -7545 5246 -7533
rect 5258 -7545 5307 -7533
rect 5187 -7637 5307 -7545
rect 5187 -7649 5247 -7637
rect 5259 -7649 5307 -7637
rect 5187 -7741 5307 -7649
rect 5187 -7753 5249 -7741
rect 5261 -7753 5307 -7741
rect 5187 -7845 5307 -7753
rect 5187 -7857 5251 -7845
rect 5263 -7857 5307 -7845
rect 5187 -7949 5307 -7857
rect 5187 -7961 5249 -7949
rect 5261 -7961 5307 -7949
rect 5187 -8053 5307 -7961
rect 5187 -8065 5246 -8053
rect 5258 -8065 5307 -8053
rect 5187 -8157 5307 -8065
rect 5187 -8169 5258 -8157
rect 5270 -8169 5307 -8157
rect 5187 -8632 5307 -8169
rect 5187 -8644 5237 -8632
rect 5249 -8644 5307 -8632
rect -3003 -13778 -111 -13096
rect 28 -13778 209 -13096
rect -3003 -13787 209 -13778
rect -3009 -14664 -663 -13998
rect -492 -14664 -323 -13998
rect -3009 -14672 -323 -14664
rect 886 -15421 1565 -15415
rect 5187 -15438 5307 -8644
rect 886 -17232 1565 -15598
rect 5304 -15752 5307 -15438
rect 5721 -7001 5841 1221
rect 9716 975 9836 985
rect 9835 659 9836 975
rect 9041 444 9161 445
rect 5721 -7089 5724 -7001
rect 5812 -7089 5841 -7001
rect 5721 -7341 5841 -7089
rect 5721 -7353 5759 -7341
rect 5771 -7353 5841 -7341
rect 5721 -7445 5841 -7353
rect 5721 -7457 5751 -7445
rect 5763 -7457 5841 -7445
rect 5721 -7549 5841 -7457
rect 5721 -7561 5742 -7549
rect 5754 -7561 5841 -7549
rect 5721 -7653 5841 -7561
rect 5721 -7665 5744 -7653
rect 5756 -7665 5841 -7653
rect 5721 -7965 5841 -7665
rect 5721 -7977 5750 -7965
rect 5762 -7977 5841 -7965
rect 5721 -8334 5841 -7977
rect 5721 -8346 5783 -8334
rect 5795 -8346 5841 -8334
rect 5721 -14758 5841 -8346
rect 6942 -103 7061 -101
rect 6942 -417 6943 -103
rect 6942 -7147 7061 -417
rect 6942 -7156 6986 -7147
rect 7009 -7156 7061 -7147
rect 6942 -14346 7061 -7156
rect 7143 -7147 7262 127
rect 8378 438 8498 442
rect 9041 128 9043 444
rect 8178 -102 8298 -101
rect 7143 -7156 7194 -7147
rect 7217 -7156 7262 -7147
rect 7143 -7666 7262 -7156
rect 8178 -7654 8298 -418
rect 7666 -7662 8298 -7654
rect 7143 -7674 7418 -7666
rect 6942 -14638 6943 -14346
rect 7143 -14758 7262 -7674
rect 8178 -14348 8298 -7662
rect 5721 -14878 7262 -14758
rect 5721 -16005 5841 -14878
rect 7143 -14899 7262 -14878
rect 8378 -14899 8498 122
rect 8841 -104 8961 -96
rect 8841 -420 8842 -104
rect 8841 -7654 8961 -420
rect 8841 -7662 8883 -7654
rect 8891 -7662 8961 -7654
rect 8841 -7726 8961 -7662
rect 8841 -7734 8863 -7726
rect 8871 -7734 8961 -7726
rect 8841 -7798 8961 -7734
rect 8841 -7806 8863 -7798
rect 8871 -7806 8961 -7798
rect 8841 -7870 8961 -7806
rect 8841 -7878 8861 -7870
rect 8869 -7878 8961 -7870
rect 8841 -7942 8961 -7878
rect 8841 -7950 8860 -7942
rect 8868 -7950 8961 -7942
rect 8841 -8014 8961 -7950
rect 8841 -8022 8861 -8014
rect 8869 -8022 8961 -8014
rect 8841 -8086 8961 -8022
rect 8841 -8094 8869 -8086
rect 8877 -8094 8961 -8086
rect 8841 -8158 8961 -8094
rect 8841 -8166 8867 -8158
rect 8875 -8166 8961 -8158
rect 8841 -14185 8961 -8166
rect 7259 -15213 7262 -14899
rect 8496 -15215 8498 -14899
rect 8378 -15221 8498 -15215
rect 8675 -14305 8961 -14185
rect 8675 -15290 8795 -14305
rect 8841 -14348 8961 -14305
rect 9041 -7594 9161 128
rect 9041 -7602 9052 -7594
rect 9060 -7602 9161 -7594
rect 9041 -7666 9161 -7602
rect 9041 -7674 9051 -7666
rect 9059 -7674 9161 -7666
rect 9041 -7738 9161 -7674
rect 9041 -7746 9061 -7738
rect 9069 -7746 9161 -7738
rect 9041 -7810 9161 -7746
rect 9041 -7818 9057 -7810
rect 9065 -7818 9161 -7810
rect 9041 -7882 9161 -7818
rect 9041 -7890 9059 -7882
rect 9067 -7890 9161 -7882
rect 9041 -7954 9161 -7890
rect 9041 -7962 9061 -7954
rect 9069 -7962 9161 -7954
rect 9041 -8026 9161 -7962
rect 9041 -8034 9060 -8026
rect 9068 -8034 9161 -8026
rect 9041 -8098 9161 -8034
rect 9041 -8106 9059 -8098
rect 9067 -8106 9161 -8098
rect 8841 -14660 8842 -14348
rect 9041 -14900 9161 -8106
rect 9716 -5502 9836 659
rect 9716 -5532 9761 -5502
rect 9791 -5532 9836 -5502
rect 9716 -5934 9836 -5532
rect 9716 -5964 9761 -5934
rect 9791 -5964 9836 -5934
rect 9716 -6370 9836 -5964
rect 9716 -6400 9761 -6370
rect 9791 -6400 9836 -6370
rect 9716 -6804 9836 -6400
rect 9716 -6834 9761 -6804
rect 9791 -6834 9836 -6804
rect 9716 -7238 9836 -6834
rect 9716 -7268 9761 -7238
rect 9791 -7268 9836 -7238
rect 9716 -7672 9836 -7268
rect 9716 -7702 9761 -7672
rect 9791 -7702 9836 -7672
rect 9716 -8106 9836 -7702
rect 9716 -8136 9761 -8106
rect 9791 -8136 9836 -8106
rect 9716 -8540 9836 -8136
rect 9716 -8570 9761 -8540
rect 9791 -8570 9836 -8540
rect 9041 -15221 9161 -15216
rect 9716 -15290 9836 -8570
rect 8675 -15410 9836 -15290
rect 9716 -15437 9836 -15410
rect 10836 -5150 10956 1224
rect 12407 973 13089 2672
rect 12407 661 13089 823
rect 14325 -1320 14510 -640
rect 14657 -1320 16677 -640
rect 13759 -2210 13945 -1533
rect 14102 -2210 16674 -1533
rect 10836 -5180 10900 -5150
rect 10930 -5180 10956 -5150
rect 10836 -5588 10956 -5180
rect 10836 -5618 10900 -5588
rect 10930 -5618 10956 -5588
rect 10836 -6017 10956 -5618
rect 10836 -6047 10901 -6017
rect 10931 -6047 10956 -6017
rect 10836 -6452 10956 -6047
rect 10836 -6482 10895 -6452
rect 10925 -6482 10956 -6452
rect 10836 -6886 10956 -6482
rect 10836 -6916 10888 -6886
rect 10918 -6916 10956 -6886
rect 10836 -7320 10956 -6916
rect 10836 -7350 10900 -7320
rect 10930 -7350 10956 -7320
rect 10836 -7754 10956 -7350
rect 10836 -7784 10894 -7754
rect 10924 -7784 10956 -7754
rect 10836 -8188 10956 -7784
rect 10836 -8218 10892 -8188
rect 10922 -8218 10956 -8188
rect 9716 -15755 9836 -15753
rect 5839 -16320 5841 -16005
rect 10836 -16007 10956 -8218
rect 14870 -13761 15035 -13086
rect 15212 -13761 16670 -13086
rect 14870 -13764 16670 -13761
rect 12444 -14532 13130 -14343
rect 12444 -14669 12447 -14532
rect 12444 -17227 13130 -14669
rect 13339 -15064 14003 -14871
rect 13339 -15230 13341 -15064
rect 13339 -17237 14003 -15230
use pad  pad_48
timestamp 1575998002
transform 1 0 -29 0 1 2000
box -3 -4 672 668
use pad  pad_49
timestamp 1575998002
transform 1 0 860 0 1 2000
box -3 -4 672 668
use pad  pad_50
timestamp 1575998002
transform 1 0 1749 0 1 2000
box -3 -4 672 668
use pad  pad_51
timestamp 1575998002
transform 1 0 2638 0 1 2000
box -3 -4 672 668
use pad  pad_52
timestamp 1575998002
transform 1 0 3527 0 1 2000
box -3 -4 672 668
use pad  pad_53
timestamp 1575998002
transform 1 0 4416 0 1 2000
box -3 -4 672 668
use pad  pad_54
timestamp 1575998002
transform 1 0 5305 0 1 2000
box -3 -4 672 668
use pad  pad_55
timestamp 1575998002
transform 1 0 6194 0 1 2000
box -3 -4 672 668
use pad  pad_56
timestamp 1575998002
transform 1 0 7083 0 1 2000
box -3 -4 672 668
use pad  pad_57
timestamp 1575998002
transform 1 0 7972 0 1 2000
box -3 -4 672 668
use pad  pad_58
timestamp 1575998002
transform 1 0 8861 0 1 2000
box -3 -4 672 668
use pad  pad_59
timestamp 1575998002
transform 1 0 9750 0 1 2000
box -3 -4 672 668
use pad  pad_60
timestamp 1575998002
transform 1 0 10639 0 1 2000
box -3 -4 672 668
use pad  pad_61
timestamp 1575998002
transform 1 0 11528 0 1 2000
box -3 -4 672 668
use pad  pad_62
timestamp 1575998002
transform 1 0 12417 0 1 2000
box -3 -4 672 668
use pad  pad_63
timestamp 1575998002
transform 1 0 13306 0 1 2000
box -3 -4 672 668
use pad  pad_32
timestamp 1575998002
transform 0 1 -2998 -1 0 -662
box -3 -4 672 668
use pad  pad_16
timestamp 1575998002
transform 0 1 16001 -1 0 -645
box -3 -4 672 668
use pad  pad_33
timestamp 1575998002
transform 0 1 -2998 -1 0 -1551
box -3 -4 672 668
use pad  pad_17
timestamp 1575998002
transform 0 1 16001 -1 0 -1534
box -3 -4 672 668
use pad  pad_34
timestamp 1575998002
transform 0 1 -2998 -1 0 -2440
box -3 -4 672 668
use pad  pad_18
timestamp 1575998002
transform 0 1 16001 -1 0 -2423
box -3 -4 672 668
use pad  pad_35
timestamp 1575998002
transform 0 1 -2998 -1 0 -3329
box -3 -4 672 668
use pad  pad_19
timestamp 1575998002
transform 0 1 16001 -1 0 -3312
box -3 -4 672 668
use pad  pad_36
timestamp 1575998002
transform 0 1 -2998 -1 0 -4218
box -3 -4 672 668
use pad  pad_20
timestamp 1575998002
transform 0 1 16001 -1 0 -4201
box -3 -4 672 668
use pad  pad_37
timestamp 1575998002
transform 0 1 -2998 -1 0 -5107
box -3 -4 672 668
use pad  pad_38
timestamp 1575998002
transform 0 1 -2998 -1 0 -5996
box -3 -4 672 668
use pad  pad_39
timestamp 1575998002
transform 0 1 -2998 -1 0 -6885
box -3 -4 672 668
use pad  pad_40
timestamp 1575998002
transform 0 1 -2998 -1 0 -7774
box -3 -4 672 668
use input_driver  input_driver_3
array 0 0 230 0 7 104
timestamp 1576130499
transform 1 0 5386 0 1 -8169
box 0 0 231 100
use input_driver  input_driver_2
array 0 0 -230 0 7 104
timestamp 1576130499
transform 0 1 6426 -1 0 -7152
box 0 0 231 100
use output_driver  output_driver_2
timestamp 1576137657
transform 0 -1 7676 1 0 -7124
box -244 -133 854 301
use core  core_0
timestamp 1576127674
transform 1 0 6186 0 1 -8168
box -322 -73 2624 656
use input_driver  input_driver_1
array 0 0 230 0 7 -104
timestamp 1576130499
transform 0 -1 6127 1 0 -8608
box 0 0 231 100
use output_driver  output_driver_0
array 0 0 1098 0 7 434
timestamp 1576137657
transform 1 0 9889 0 1 -8454
box -244 -133 854 301
use pad  pad_21
timestamp 1575998002
transform 0 1 16001 -1 0 -5090
box -3 -4 672 668
use pad  pad_22
timestamp 1575998002
transform 0 1 16001 -1 0 -5979
box -3 -4 672 668
use pad  pad_23
timestamp 1575998002
transform 0 1 16001 -1 0 -6868
box -3 -4 672 668
use pad  pad_24
timestamp 1575998002
transform 0 1 16001 -1 0 -7757
box -3 -4 672 668
use pad  pad_41
timestamp 1575998002
transform 0 1 -2998 -1 0 -8663
box -3 -4 672 668
use pad  pad_42
timestamp 1575998002
transform 0 1 -2998 -1 0 -9552
box -3 -4 672 668
use output_driver  output_driver_1
array 0 0 -1098 0 6 434
timestamp 1576137657
transform 0 1 7046 -1 0 -8902
box -244 -133 854 301
use pad  pad_25
timestamp 1575998002
transform 0 1 16001 -1 0 -8646
box -3 -4 672 668
use pad  pad_26
timestamp 1575998002
transform 0 1 16001 -1 0 -9535
box -3 -4 672 668
use pad  pad_43
timestamp 1575998002
transform 0 1 -2998 -1 0 -10441
box -3 -4 672 668
use pad  pad_27
timestamp 1575998002
transform 0 1 16001 -1 0 -10424
box -3 -4 672 668
use pad  pad_44
timestamp 1575998002
transform 0 1 -2998 -1 0 -11330
box -3 -4 672 668
use pad  pad_28
timestamp 1575998002
transform 0 1 16001 -1 0 -11313
box -3 -4 672 668
use pad  pad_45
timestamp 1575998002
transform 0 1 -2998 -1 0 -12219
box -3 -4 672 668
use pad  pad_29
timestamp 1575998002
transform 0 1 16001 -1 0 -12202
box -3 -4 672 668
use pad  pad_46
timestamp 1575998002
transform 0 1 -2998 -1 0 -13108
box -3 -4 672 668
use pad  pad_30
timestamp 1575998002
transform 0 1 16001 -1 0 -13091
box -3 -4 672 668
use pad  pad_47
timestamp 1575998002
transform 0 1 -2998 -1 0 -13997
box -3 -4 672 668
use pad  pad_31
timestamp 1575998002
transform 0 1 16001 -1 0 -13980
box -3 -4 672 668
use pad  pad_0
timestamp 1575998002
transform 1 0 0 0 1 -17223
box -3 -4 672 668
use pad  pad_1
timestamp 1575998002
transform 1 0 889 0 1 -17223
box -3 -4 672 668
use pad  pad_2
timestamp 1575998002
transform 1 0 1778 0 1 -17223
box -3 -4 672 668
use pad  pad_3
timestamp 1575998002
transform 1 0 2667 0 1 -17223
box -3 -4 672 668
use pad  pad_4
timestamp 1575998002
transform 1 0 3556 0 1 -17223
box -3 -4 672 668
use pad  pad_5
timestamp 1575998002
transform 1 0 4445 0 1 -17223
box -3 -4 672 668
use pad  pad_6
timestamp 1575998002
transform 1 0 5334 0 1 -17223
box -3 -4 672 668
use pad  pad_7
timestamp 1575998002
transform 1 0 6223 0 1 -17223
box -3 -4 672 668
use pad  pad_8
timestamp 1575998002
transform 1 0 7112 0 1 -17223
box -3 -4 672 668
use pad  pad_9
timestamp 1575998002
transform 1 0 8001 0 1 -17223
box -3 -4 672 668
use pad  pad_10
timestamp 1575998002
transform 1 0 8890 0 1 -17223
box -3 -4 672 668
use pad  pad_11
timestamp 1575998002
transform 1 0 9779 0 1 -17223
box -3 -4 672 668
use pad  pad_12
timestamp 1575998002
transform 1 0 10668 0 1 -17223
box -3 -4 672 668
use pad  pad_13
timestamp 1575998002
transform 1 0 11557 0 1 -17223
box -3 -4 672 668
use pad  pad_14
timestamp 1575998002
transform 1 0 12446 0 1 -17223
box -3 -4 672 668
use pad  pad_15
timestamp 1575998002
transform 1 0 13335 0 1 -17223
box -3 -4 672 668
<< labels >>
rlabel metal5 10829 -5360 10829 -5360 1 d0
rlabel metal5 10829 -5787 10829 -5787 1 d1
rlabel metal5 10820 -6236 10820 -6236 1 d2
rlabel metal5 10818 -6643 10818 -6643 1 d3
rlabel metal5 10811 -7097 10811 -7097 1 d4
rlabel metal5 10811 -7541 10811 -7541 1 d5
rlabel metal5 10805 -7983 10805 -7983 1 d6
rlabel metal5 10795 -8400 10795 -8400 1 d7
rlabel m4contact 9342 -9768 9342 -9768 1 c6
rlabel m4contact 8007 -9771 8007 -9771 1 c3
rlabel m4contact 7588 -9768 7588 -9768 1 c2
rlabel m4contact 7142 -9767 7142 -9767 1 c1
rlabel m4contact 6804 -8613 6804 -8613 1 b7
rlabel m4contact 6701 -8612 6701 -8612 1 b6
rlabel m4contact 6594 -8612 6594 -8612 1 opcode2
rlabel m4contact 6490 -8610 6490 -8610 1 b5
rlabel m4contact 6386 -8611 6386 -8611 1 Den
rlabel m4contact 6283 -8610 6283 -8610 1 opcode1
rlabel m4contact 6179 -8612 6179 -8612 1 Cen
rlabel m4contact 6076 -8611 6076 -8611 1 opcode0
rlabel m4contact 5380 -8118 5380 -8118 1 clk
rlabel m4contact 5382 -8014 5382 -8014 1 Bctrl
rlabel m4contact 5381 -7910 5381 -7910 1 Actrl
rlabel m4contact 5380 -7806 5380 -7806 1 b4
rlabel m4contact 5380 -7701 5380 -7701 1 b3
rlabel m4contact 5380 -7598 5380 -7598 1 b2
rlabel m4contact 5380 -7493 5380 -7493 1 b1
rlabel m4contact 5378 -7391 5378 -7391 1 b0
rlabel m4contact 9690 -9766 9690 -9766 1 c7
rlabel m4contact 8824 -9766 8824 -9766 1 c5
rlabel m4contact 8511 -9770 8511 -9770 1 c4
rlabel metal4 6456 -7148 6456 -7148 1 a0
rlabel m4contact 6582 -7151 6582 -7151 1 a1
rlabel m4contact 6686 -7151 6687 -7151 1 a2
rlabel m4contact 6788 -7151 6788 -7151 1 a3
rlabel m4contact 6893 -7150 6893 -7150 1 a4
rlabel m4contact 6997 -7151 6997 -7151 1 a5
rlabel m4contact 7100 -7151 7100 -7151 1 a6
rlabel m4contact 7205 -7151 7205 -7151 1 a7
rlabel metal4 7687 -14502 7687 -14502 1 Gnd
rlabel metal4 7665 -15059 7665 -15059 1 Vdd
rlabel metal4 7643 -15599 7643 -15599 1 Gnd
rlabel metal4 7632 -16182 7632 -16182 1 Vdd
rlabel m345contact 7597 -6268 7597 -6268 1 c0
rlabel m4contact 7094 -7389 7094 -7389 1 _a6
rlabel m4contact 6186 -8368 6186 -8368 1 _cen
rlabel metal5 8650 -8155 8650 -8155 1 nz7
rlabel metal5 8813 -8148 8813 -8148 1 _d7
rlabel metal1 10102 -8427 10102 -8427 1 _drv_d7
<< end >>
