magic
tech scmos
timestamp 1575778961
<< error_s >>
rect 308 445 318 446
rect 548 373 558 374
rect 788 301 798 302
rect 1028 229 1038 230
rect 1268 157 1278 158
rect 1508 85 1518 86
rect 1748 13 1758 14
<< m4contact >>
rect -117 463 -108 472
rect 123 391 132 400
rect 363 318 372 327
rect 603 246 612 255
rect 843 174 852 183
rect 1083 102 1092 111
rect 1143 31 1152 40
rect 1323 31 1332 40
<< metal4 >>
rect -117 472 -108 553
rect 123 400 132 481
rect 363 327 372 409
rect 603 255 612 337
rect 843 183 852 265
rect 1083 111 1092 193
rect 1143 40 1152 121
rect 1323 40 1332 49
<< m5contact >>
rect -117 553 -108 562
rect 123 481 132 490
rect 363 409 372 418
rect 603 337 612 346
rect 843 265 852 274
rect 1083 193 1092 202
rect 1143 121 1152 130
rect 1323 49 1332 58
<< metal6 >>
rect 1874 62 1882 593
rect 1890 2 1898 593
use logic  logic_0
timestamp 1575777673
transform 1 0 -327 0 1 504
box 87 2 327 70
use fadder  fadder_0
timestamp 1575778664
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1575777673
transform 1 0 -87 0 1 432
box 87 2 327 70
use fadder  fadder_1
timestamp 1575778664
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1575777673
transform 1 0 153 0 1 360
box 87 2 327 70
use fadder  fadder_2
timestamp 1575778664
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1575777673
transform 1 0 393 0 1 288
box 87 2 327 70
use fadder  fadder_3
timestamp 1575778664
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1575777673
transform 1 0 633 0 1 216
box 87 2 327 70
use fadder  fadder_4
timestamp 1575778664
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1575777673
transform 1 0 873 0 1 144
box 87 2 327 70
use fadder  fadder_5
timestamp 1575778664
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1575777673
transform 1 0 1113 0 1 72
box 87 2 327 70
use fadder  fadder_6
timestamp 1575778664
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1575778664
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1575777673
transform 1 0 1353 0 1 0
box 87 2 327 70
use mult  mult_0
timestamp 1575778961
transform 1 0 241 0 1 432
box -481 -432 1679 142
<< labels >>
rlabel metal6 1878 590 1878 590 5 Vdd
rlabel metal6 1894 589 1894 589 5 Gnd
<< end >>
