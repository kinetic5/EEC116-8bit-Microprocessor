magic
tech scmos
timestamp 1575941385
<< ntransistor >>
rect -19 21 -17 27
rect -9 23 -7 27
rect -29 12 -27 16
<< ptransistor >>
rect -29 50 -27 56
rect -19 39 -17 45
rect -9 39 -7 45
<< ndiffusion >>
rect -26 25 -19 27
rect -26 21 -25 25
rect -20 21 -19 25
rect -17 23 -15 27
rect -10 23 -9 27
rect -7 23 -6 27
rect -17 21 -13 23
rect -31 15 -29 16
rect -36 12 -29 15
rect -27 12 -21 16
rect -26 8 -21 12
<< pdiffusion >>
rect -26 56 -21 60
rect -30 50 -29 56
rect -27 50 -21 56
rect -20 40 -19 45
rect -26 39 -19 40
rect -17 39 -15 45
rect -10 39 -9 45
rect -7 39 -6 45
<< ndcontact >>
rect -36 15 -31 19
rect -25 21 -20 25
rect -15 23 -10 27
rect -26 4 -21 8
<< pdcontact >>
rect -26 60 -20 64
rect -36 50 -30 56
rect -26 40 -20 45
rect -15 39 -10 45
<< polysilicon >>
rect -39 11 -37 57
rect -29 56 -27 59
rect -19 53 -17 57
rect -9 54 -7 57
rect -29 32 -27 50
rect -19 45 -17 48
rect -9 45 -7 49
rect -19 36 -17 39
rect -9 36 -7 39
rect -29 16 -27 28
rect -19 27 -17 30
rect -9 27 -7 30
rect -19 18 -17 21
rect -9 17 -7 23
rect -29 9 -27 12
rect -19 11 -17 13
rect -9 11 -7 12
<< polycontact >>
rect -31 28 -27 32
<< metal1 >>
rect -43 64 -3 68
rect -43 60 -26 64
rect -20 60 -3 64
rect -41 50 -36 56
rect -30 50 -29 56
rect -41 26 -35 50
rect -20 40 -18 45
rect -36 21 -35 26
rect -20 21 -18 25
rect -15 35 -10 39
rect -15 30 8 35
rect -15 27 -10 30
rect -41 19 -35 21
rect -41 15 -36 19
rect -43 4 -26 8
rect -21 4 -1 8
rect -43 0 -1 4
<< pm12contact >>
rect -20 48 -15 53
rect -11 49 -6 54
rect -20 13 -15 18
rect -11 12 -6 17
<< pdm12contact >>
rect -6 39 0 45
<< ndm12contact >>
rect -6 21 0 27
<< metal2 >>
rect -41 48 -20 53
rect -41 26 -36 48
rect -32 18 -27 32
rect -32 13 -20 18
<< m3contact >>
rect -6 49 -1 54
rect -6 27 0 39
rect -6 12 -1 17
<< m123contact >>
rect -41 21 -36 26
rect -32 32 -27 37
rect -23 25 -18 40
<< metal3 >>
rect -32 49 -6 54
rect -32 37 -27 49
rect 92 40 100 48
rect -41 17 -36 21
rect -41 12 -6 17
use dff  dff_0
timestamp 1575941385
transform 1 0 -3 0 1 61
box 0 -61 150 7
<< labels >>
rlabel m3contact -3 33 -3 33 1 in_0
rlabel m123contact -21 32 -21 32 1 in_1
rlabel m123contact -30 34 -30 34 1 enable
rlabel metal1 -15 4 -15 4 1 Gnd
rlabel metal1 -14 64 -14 64 5 Vdd
rlabel metal1 -13 32 -13 32 1 mux_out
rlabel metal3 96 47 96 47 1 clk
<< end >>
