magic
tech scmos
timestamp 1576132548
<< nwell >>
rect 136 29 195 68
<< pwell >>
rect 419 140 435 161
rect 136 -4 200 29
<< ntransistor >>
rect 150 13 152 23
rect 160 13 162 23
rect 170 13 172 23
rect 180 13 182 23
<< ptransistor >>
rect 150 37 152 51
rect 160 37 162 51
rect 170 37 172 51
rect 180 37 182 51
<< ndiffusion >>
rect 149 13 150 23
rect 152 22 160 23
rect 152 13 153 22
rect 159 13 160 22
rect 162 13 163 23
rect 169 13 170 23
rect 172 13 173 23
rect 179 13 180 23
rect 182 13 183 23
rect 189 11 190 23
<< pdiffusion >>
rect 149 37 150 51
rect 152 38 153 51
rect 159 38 160 51
rect 152 37 160 38
rect 162 37 163 51
rect 169 37 170 51
rect 172 37 173 51
rect 179 37 180 51
rect 182 37 183 51
<< ndcontact >>
rect 143 13 149 23
rect 163 13 169 23
rect 183 11 189 23
<< pdcontact >>
rect 143 37 149 51
rect 163 37 169 51
rect 183 35 189 53
<< psubstratepcontact >>
rect 140 -1 152 6
rect 171 -1 183 6
<< nsubstratencontact >>
rect 140 58 152 65
rect 171 58 183 65
<< polysilicon >>
rect 140 8 142 56
rect 150 51 152 56
rect 160 51 162 56
rect 170 51 172 56
rect 180 51 182 56
rect 150 32 152 37
rect 160 32 162 37
rect 170 32 172 37
rect 180 32 182 37
rect 150 23 152 26
rect 160 23 162 26
rect 170 23 172 26
rect 180 23 182 26
rect 150 8 152 13
rect 160 8 162 13
rect 170 8 172 13
rect 180 8 182 13
<< polycontact >>
rect 158 26 164 32
rect 168 26 174 32
rect 178 26 184 32
<< metal1 >>
rect 136 65 193 66
rect 136 58 140 65
rect 152 58 171 65
rect 183 58 193 65
rect 143 51 149 58
rect 163 51 169 58
rect 183 53 189 58
rect 147 26 148 32
rect 154 26 158 32
rect 164 26 168 32
rect 174 26 178 32
rect 143 6 149 13
rect 163 6 169 13
rect 183 6 189 11
rect 136 -1 140 6
rect 152 -1 171 6
rect 183 -1 193 6
rect 136 -2 193 -1
<< pm12contact >>
rect 148 26 154 32
<< pdm12contact >>
rect 153 38 159 51
rect 173 37 179 51
<< ndm12contact >>
rect 153 13 159 22
rect 173 13 179 23
<< metal2 >>
rect 166 62 175 68
rect 159 37 173 51
rect 179 49 183 51
rect 179 45 189 49
rect 142 32 148 33
rect 147 26 148 32
rect 142 25 148 26
rect 179 25 189 35
rect 159 13 173 23
rect 179 13 189 15
rect 165 -4 174 2
<< m3contact >>
rect 142 33 148 38
rect 179 35 189 45
rect 142 20 148 25
rect 179 15 189 25
<< m123contact >>
rect 142 26 147 32
<< metal3 >>
rect 142 32 148 33
rect 147 26 148 32
rect 142 25 148 26
rect 179 25 189 35
<< end >>
