magic
tech scmos
timestamp 1576006893
<< nwell >>
rect 13 101 232 244
<< pwell >>
rect 13 -77 231 47
<< ntransistor >>
rect 47 -20 49 20
rect 57 -20 59 20
rect 67 -20 69 20
rect 77 -20 79 20
rect 87 -20 89 20
rect 97 -20 99 20
rect 107 -20 109 20
rect 117 -20 119 20
rect 127 -20 129 20
rect 137 -20 139 20
rect 147 -20 149 20
rect 157 -20 159 20
rect 167 -20 169 20
rect 177 -20 179 20
rect 187 -20 189 20
rect 197 -20 199 20
<< ptransistor >>
rect 47 132 49 192
rect 57 132 59 192
rect 67 132 69 192
rect 77 132 79 192
rect 87 132 89 192
rect 97 132 99 192
rect 107 132 109 192
rect 117 132 119 192
rect 127 132 129 192
rect 137 132 139 192
rect 147 132 149 192
rect 157 132 159 192
rect 167 132 169 192
rect 177 132 179 192
rect 187 132 189 192
rect 197 132 199 192
<< ndiffusion >>
rect 46 -20 47 20
rect 49 -20 50 20
rect 56 -20 57 20
rect 59 -20 60 20
rect 66 -20 67 20
rect 69 -20 70 20
rect 76 -20 77 20
rect 79 -20 80 20
rect 86 -20 87 20
rect 89 -20 90 20
rect 96 -20 97 20
rect 99 -20 100 20
rect 106 -20 107 20
rect 109 -20 110 20
rect 116 -20 117 20
rect 119 -20 120 20
rect 126 -20 127 20
rect 129 -20 130 20
rect 136 -20 137 20
rect 139 -20 140 20
rect 146 -20 147 20
rect 149 -20 150 20
rect 156 -20 157 20
rect 159 -20 160 20
rect 166 -20 167 20
rect 169 -20 170 20
rect 176 -20 177 20
rect 179 -20 180 20
rect 186 -20 187 20
rect 189 -20 190 20
rect 196 -20 197 20
rect 199 -20 200 20
<< pdiffusion >>
rect 46 132 47 192
rect 49 132 50 192
rect 56 132 57 192
rect 59 132 60 192
rect 66 132 67 192
rect 69 132 70 192
rect 76 132 77 192
rect 79 132 80 192
rect 86 132 87 192
rect 89 132 90 192
rect 96 132 97 192
rect 99 132 100 192
rect 106 132 107 192
rect 109 132 110 192
rect 116 132 117 192
rect 119 132 120 192
rect 126 132 127 192
rect 129 132 130 192
rect 136 132 137 192
rect 139 132 140 192
rect 146 132 147 192
rect 149 132 150 192
rect 156 132 157 192
rect 159 132 160 192
rect 166 132 167 192
rect 169 132 170 192
rect 176 132 177 192
rect 179 132 180 192
rect 186 132 187 192
rect 189 132 190 192
rect 196 132 197 192
rect 199 132 200 192
<< ndcontact >>
rect 40 -20 46 20
rect 60 -20 66 20
rect 80 -20 86 20
rect 100 -20 106 20
rect 120 -20 126 20
rect 140 -20 146 20
rect 160 -20 166 20
rect 180 -20 186 20
rect 200 -20 206 20
<< pdcontact >>
rect 40 132 46 192
rect 60 132 66 192
rect 80 132 86 192
rect 100 132 106 192
rect 120 132 126 192
rect 140 132 146 192
rect 160 132 166 192
rect 180 132 186 192
rect 200 132 206 192
<< psubstratepcontact >>
rect 26 -52 62 -33
rect 94 -52 130 -33
rect 158 -52 194 -33
<< nsubstratencontact >>
rect 24 204 61 223
rect 99 204 136 223
rect 159 204 196 223
<< polysilicon >>
rect 47 192 49 199
rect 57 192 59 199
rect 67 192 69 199
rect 77 192 79 199
rect 87 192 89 199
rect 97 192 99 199
rect 107 192 109 199
rect 117 192 119 199
rect 127 192 129 199
rect 137 192 139 199
rect 147 192 149 199
rect 157 192 159 199
rect 167 192 169 199
rect 177 192 179 199
rect 187 192 189 199
rect 197 192 199 199
rect 47 119 49 132
rect 57 119 59 132
rect 67 119 69 132
rect 77 119 79 132
rect 87 119 89 132
rect 97 119 99 132
rect 107 119 109 132
rect 117 119 119 132
rect 127 119 129 132
rect 137 119 139 132
rect 147 119 149 132
rect 157 119 159 132
rect 167 119 169 132
rect 177 119 179 132
rect 187 119 189 132
rect 197 119 199 132
rect 47 20 49 30
rect 57 20 59 30
rect 67 20 69 30
rect 77 20 79 30
rect 87 20 89 30
rect 97 20 99 30
rect 107 20 109 30
rect 117 20 119 30
rect 127 20 129 30
rect 137 20 139 30
rect 147 20 149 30
rect 157 20 159 30
rect 167 20 169 30
rect 177 20 179 30
rect 187 20 189 30
rect 197 20 199 30
rect 47 -27 49 -20
rect 57 -27 59 -20
rect 67 -27 69 -20
rect 77 -27 79 -20
rect 87 -27 89 -20
rect 97 -27 99 -20
rect 107 -27 109 -20
rect 117 -27 119 -20
rect 127 -27 129 -20
rect 137 -27 139 -20
rect 147 -27 149 -20
rect 157 -27 159 -20
rect 167 -27 169 -20
rect 177 -27 179 -20
rect 187 -27 189 -20
rect 197 -27 199 -20
<< polycontact >>
rect 45 30 51 119
rect 55 30 61 119
rect 65 30 71 119
rect 75 30 81 119
rect 85 30 91 119
rect 95 30 101 119
rect 105 30 111 119
rect 115 30 121 119
rect 125 30 131 119
rect 135 30 141 119
rect 145 30 151 119
rect 155 30 161 119
rect 165 30 171 119
rect 175 30 181 119
rect 185 30 191 119
rect 195 30 201 119
<< metal1 >>
rect -40 223 221 227
rect -40 204 24 223
rect 61 204 99 223
rect 136 204 159 223
rect 196 204 221 223
rect -40 200 221 204
rect -40 123 -13 200
rect 40 192 46 200
rect 60 192 66 200
rect 80 192 86 200
rect 100 192 106 200
rect 120 192 126 200
rect 140 192 146 200
rect 160 192 166 200
rect 180 192 186 200
rect 200 192 206 200
rect -41 -29 -14 47
rect 2 30 45 119
rect 51 30 55 119
rect 61 30 65 119
rect 71 30 75 119
rect 81 30 85 119
rect 91 30 95 119
rect 101 30 105 119
rect 111 30 115 119
rect 121 30 125 119
rect 131 30 135 119
rect 141 30 145 119
rect 151 30 155 119
rect 161 30 165 119
rect 171 30 175 119
rect 181 30 185 119
rect 191 30 195 119
rect 201 30 202 119
rect 40 -29 46 -20
rect 60 -29 66 -20
rect 80 -29 86 -20
rect 100 -29 106 -20
rect 120 -29 126 -20
rect 140 -29 146 -20
rect 160 -29 166 -20
rect 180 -29 186 -20
rect 200 -29 206 -20
rect -41 -33 214 -29
rect -41 -52 26 -33
rect 62 -52 94 -33
rect 130 -52 158 -33
rect 194 -52 214 -33
rect -41 -56 214 -52
<< pdm12contact >>
rect 50 132 56 192
rect 70 132 76 192
rect 90 132 96 192
rect 110 132 116 192
rect 130 132 136 192
rect 150 132 156 192
rect 170 132 176 192
rect 190 132 196 192
<< ndm12contact >>
rect 50 -20 56 20
rect 70 -20 76 20
rect 90 -20 96 20
rect 110 -20 116 20
rect 130 -20 136 20
rect 150 -20 156 20
rect 170 -20 176 20
rect 190 -20 196 20
<< metal2 >>
rect 56 132 70 192
rect 76 132 90 192
rect 96 132 110 192
rect 116 132 130 192
rect 136 132 150 192
rect 156 132 170 192
rect 176 132 190 192
rect 196 132 228 192
rect -37 52 -28 118
rect 50 20 228 132
rect 56 -20 70 20
rect 76 -20 90 20
rect 96 -20 110 20
rect 116 -20 130 20
rect 136 -20 150 20
rect 156 -20 170 20
rect 176 -20 190 20
rect 196 -20 228 20
<< m3contact >>
rect 228 30 273 119
<< m123contact >>
rect -12 52 2 118
<< metal3 >>
rect -30 52 -12 118
use input_driver  input_driver_0
timestamp 1576001165
transform 1 0 -244 0 1 35
box 0 0 230 100
<< labels >>
rlabel m3contact 267 71 267 71 1 out
<< end >>
