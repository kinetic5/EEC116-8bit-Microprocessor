magic
tech scmos
timestamp 1576125678
<< error_p >>
rect 6564 -7175 6565 -7169
rect 6564 -7195 6565 -7189
rect 6564 -7215 6565 -7209
rect 6564 -7265 6565 -7219
rect 5403 -8031 5409 -8030
rect 5423 -8031 5429 -8030
rect 5443 -8031 5449 -8030
rect 5453 -8031 5499 -8030
rect 9912 -8172 9913 -8171
rect 9911 -8173 9912 -8172
rect 9915 -8191 9916 -8190
rect 9914 -8192 9915 -8191
rect 6092 -8541 6093 -8495
rect 6092 -8551 6093 -8545
rect 6092 -8571 6093 -8565
rect 6092 -8591 6093 -8585
<< error_s >>
rect 6876 -7175 6877 -7169
rect 6980 -7175 6981 -7169
rect 7084 -7175 7085 -7169
rect 7188 -7175 7189 -7169
rect 6876 -7195 6877 -7189
rect 6980 -7195 6981 -7189
rect 7084 -7195 7085 -7189
rect 7188 -7195 7189 -7189
rect 6876 -7215 6877 -7209
rect 6980 -7215 6981 -7209
rect 7084 -7215 7085 -7209
rect 7188 -7215 7189 -7209
rect 6876 -7265 6877 -7219
rect 6980 -7265 6981 -7219
rect 7084 -7265 7085 -7219
rect 7188 -7265 7189 -7219
rect 8405 -7710 8406 -7709
rect 8405 -7783 8406 -7779
rect 5865 -7841 5866 -7840
rect 5866 -7849 5867 -7841
rect 5865 -7850 5866 -7849
rect 8796 -7910 8804 -7909
rect 8797 -7984 8805 -7981
rect 6196 -8541 6197 -8495
rect 6300 -8541 6301 -8495
rect 6820 -8541 6821 -8495
rect 6196 -8551 6197 -8545
rect 6300 -8551 6301 -8545
rect 6820 -8551 6821 -8545
rect 6196 -8571 6197 -8565
rect 6300 -8571 6301 -8565
rect 6820 -8571 6821 -8565
rect 6196 -8591 6197 -8585
rect 6300 -8591 6301 -8585
rect 6820 -8591 6821 -8585
rect 8195 -8925 8196 -8924
rect 9063 -8925 9064 -8924
rect 8196 -8926 8197 -8925
rect 9064 -8926 9065 -8925
rect 8176 -8928 8177 -8927
rect 9044 -8928 9045 -8927
rect 8177 -8929 8178 -8928
rect 9045 -8929 9046 -8928
<< error_ps >>
rect 7327 -8925 7328 -8924
rect 7328 -8926 7329 -8925
rect 7308 -8928 7309 -8927
rect 7309 -8929 7310 -8928
<< pwell >>
rect 6083 -8508 6125 -8485
rect 6083 -8527 6087 -8508
rect 6083 -8608 6125 -8527
<< metal1 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1543 13975 1569
rect -1773 1541 15766 1543
rect -1773 1529 15098 1541
rect -1773 1232 -1767 1529
rect -754 1232 15098 1529
rect -1773 1214 15098 1232
rect -1773 226 -1444 1214
rect 15425 1214 15766 1541
rect 15437 1197 15766 1214
rect -1773 -623 -1772 226
rect -1449 -623 -1444 226
rect -1773 -654 -1444 -623
rect -1216 657 14878 986
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -1336 -1441 -665
rect -3013 -1341 -1441 -1336
rect -1773 -15993 -1444 -1341
rect -1216 -15423 -887 657
rect 232 650 561 657
rect 14873 645 14878 657
rect 15437 868 15441 1197
rect 232 456 561 457
rect -667 127 14661 456
rect -666 -14873 -337 127
rect -116 -95 213 -94
rect 577 -95 14100 -94
rect -116 -423 14100 -95
rect -116 -14336 213 -423
rect 13771 -3679 14100 -423
rect 13756 -4525 14100 -3679
rect 8810 -7602 9068 -7594
rect 8810 -7662 8899 -7654
rect 8810 -7674 9067 -7666
rect 9075 -7674 9076 -7666
rect 8810 -7734 8879 -7726
rect 8887 -7734 8927 -7726
rect 8810 -7746 9077 -7738
rect 8810 -7806 8879 -7798
rect 8810 -7818 9073 -7810
rect 8810 -7878 8877 -7870
rect 8810 -7890 9075 -7882
rect 8810 -7950 8876 -7942
rect 8809 -7962 9077 -7954
rect 8810 -8022 8877 -8014
rect 8810 -8034 9076 -8026
rect 8810 -8094 8885 -8086
rect 8810 -8106 9075 -8098
rect 8810 -8166 8883 -8158
rect 13756 -14333 14085 -4525
rect -116 -14341 222 -14336
rect 582 -14341 13655 -14336
rect -116 -14658 13655 -14341
rect -116 -14665 222 -14658
rect 588 -14665 13655 -14658
rect 14323 -14871 14655 127
rect 14873 -1424 15202 645
rect 232 -14873 561 -14872
rect 866 -14873 14655 -14871
rect -666 -14876 14655 -14873
rect -666 -15202 14211 -14876
rect -664 -15211 14211 -15202
rect 14645 -15200 14655 -14876
rect 14870 -3055 15202 -1424
rect 14870 -14709 15199 -3055
rect 15437 -13974 15766 868
rect 15434 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 14870 -15053 14871 -14709
rect 15437 -14766 15766 -14654
rect 14645 -15211 14649 -15200
rect 14870 -15418 15199 -15053
rect 232 -15423 561 -15420
rect -1216 -15752 14778 -15423
rect 15521 -14799 15766 -14766
rect 15521 -15983 15646 -14799
rect 15437 -15989 15646 -15983
rect 10 -15993 661 -15992
rect 15437 -15993 15768 -15989
rect -1773 -15998 8414 -15993
rect -1773 -16081 14470 -15998
rect -1773 -16210 15766 -16081
rect -1773 -16315 14469 -16210
rect -1773 -16322 10 -16315
rect 661 -16322 14469 -16315
rect 7835 -16324 14469 -16322
rect 15753 -16324 15766 -16210
rect 7835 -16327 15766 -16324
rect 10 -17229 661 -16553
<< metal2 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1546 13975 1569
rect 240 1543 15763 1546
rect -1774 1541 15763 1543
rect -1774 1538 15098 1541
rect -1774 1529 13299 1538
rect -1774 1232 -1767 1529
rect -754 1232 13299 1529
rect -1774 1217 13299 1232
rect -1774 1214 890 1217
rect -1774 1211 -1445 1214
rect -1774 255 -1767 1211
rect -1456 255 -1445 1211
rect 13971 1217 15098 1538
rect 15425 1219 15436 1541
rect 15758 1219 15763 1541
rect 15425 1217 15763 1219
rect 15434 1197 15763 1217
rect -929 981 14512 982
rect -1774 226 -1445 255
rect -1774 -623 -1772 226
rect -1449 -623 -1445 226
rect -1774 -654 -1445 -623
rect -1217 814 14512 981
rect -1217 664 12407 814
rect 13092 664 14512 814
rect -1217 660 14512 664
rect 14852 660 14878 982
rect -1217 653 14878 660
rect -1217 652 896 653
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -670 -1441 -665
rect -1835 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -1835 -1336 -1441 -1331
rect -3013 -1341 -1441 -1336
rect -1774 -15992 -1445 -1341
rect -1217 -1544 -888 652
rect 15434 868 15441 1197
rect 14884 618 15213 645
rect -1217 -2224 -1047 -1544
rect -889 -2224 -888 -1544
rect -1217 -15428 -888 -2224
rect -667 444 876 457
rect -667 129 14649 444
rect -667 -14001 -339 129
rect 467 116 14649 129
rect 1720 -95 2049 -94
rect 2520 -95 14096 -93
rect -116 -422 14096 -95
rect -116 -423 3442 -422
rect -116 -424 222 -423
rect 582 -424 3442 -423
rect -116 -13100 213 -424
rect 13767 -1532 14096 -422
rect 13932 -2213 14096 -1532
rect -116 -13787 42 -13100
rect 200 -13787 213 -13100
rect -667 -14674 -482 -14001
rect -116 -14333 213 -13787
rect 13767 -13979 14096 -2213
rect 14095 -14312 14096 -13979
rect 13767 -14333 14096 -14312
rect 14321 -636 14649 116
rect 14321 -1321 14327 -636
rect 14499 -1321 14649 -636
rect -116 -14341 222 -14333
rect 582 -14341 13267 -14333
rect -116 -14347 13267 -14341
rect -116 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -116 -14662 13267 -14484
rect 13646 -14662 13655 -14333
rect 14321 -14517 14649 -1321
rect 14884 -13082 15213 272
rect 15028 -13769 15213 -13082
rect -667 -14883 -339 -14674
rect 14321 -14850 14327 -14517
rect 14884 -14709 15213 -13769
rect 14321 -14876 14649 -14850
rect -667 -15043 13336 -14883
rect 14002 -15043 14211 -14883
rect -667 -15211 14211 -15043
rect 14645 -15211 14649 -14876
rect 15212 -15053 15213 -14709
rect 14884 -15063 15213 -15053
rect 15212 -15398 15213 -15063
rect 14884 -15418 15213 -15398
rect -1217 -15609 14338 -15428
rect -1217 -15757 886 -15609
rect 1567 -15757 14338 -15609
rect 14772 -15757 14778 -15428
rect 15212 -15757 15213 -15418
rect 15434 -13972 15763 868
rect 15434 -14674 15436 -13972
rect 15747 -13974 15763 -13972
rect 15747 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 15747 -14674 15763 -14654
rect 15434 -14694 15763 -14674
rect 15434 -14766 15766 -14694
rect 15521 -14771 15766 -14766
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -14799 15766 -14771
rect 15644 -15986 15646 -14799
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16081 14470 -15993
rect 662 -16090 15766 -16081
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16210 15766 -16204
rect 662 -16313 14469 -16210
rect -1774 -16315 14469 -16313
rect -1774 -16321 10 -16315
rect -9 -16322 10 -16321
rect 661 -16321 14469 -16315
rect 15753 -16321 15766 -16210
rect 10 -17229 661 -16553
<< m123contact >>
rect 13308 1569 13962 1943
rect -1767 1232 -754 1529
rect 15098 1212 15425 1541
rect -1772 -623 -1449 226
rect -2255 -1336 -1835 -665
rect 14878 645 15219 991
rect 15441 868 15768 1197
rect 8488 -7602 8496 -7594
rect 9068 -7602 9076 -7594
rect 7642 -7660 7650 -7654
rect 8899 -7662 8907 -7654
rect 7402 -7672 7410 -7666
rect 8487 -7674 8495 -7668
rect 9067 -7674 9075 -7666
rect 8879 -7734 8887 -7726
rect 9077 -7746 9085 -7738
rect 7591 -7804 7599 -7798
rect 8628 -7804 8636 -7798
rect 8879 -7806 8887 -7798
rect 9073 -7818 9081 -7810
rect 8632 -7876 8640 -7870
rect 8877 -7878 8885 -7870
rect 8686 -7888 8694 -7882
rect 9075 -7890 9083 -7882
rect 8647 -7948 8655 -7942
rect 8876 -7950 8884 -7942
rect 8683 -7960 8691 -7954
rect 9077 -7962 9085 -7954
rect 8632 -8020 8640 -8014
rect 8877 -8022 8885 -8014
rect 9076 -8034 9084 -8026
rect 8681 -8092 8689 -8086
rect 8885 -8094 8893 -8086
rect 8638 -8104 8646 -8098
rect 9075 -8106 9083 -8098
rect 8655 -8164 8663 -8158
rect 8883 -8166 8891 -8158
rect 13655 -14672 14099 -14333
rect 14211 -15222 14645 -14876
rect 14871 -15053 15212 -14709
rect 14778 -15764 15212 -15418
rect 15766 -14654 15975 -13974
rect 15434 -15983 15521 -14766
rect 15646 -15989 15768 -14799
rect 14470 -16081 15768 -15993
rect 10 -16553 661 -16315
rect 14469 -16324 15753 -16210
<< metal3 >>
rect 13304 1943 13975 2669
rect 13304 1569 13308 1943
rect 13962 1569 13975 1943
rect 13304 1546 13975 1569
rect -1774 1541 15763 1546
rect -1774 1538 15098 1541
rect -1774 1529 13299 1538
rect -1774 1232 -1767 1529
rect -754 1232 13299 1529
rect -1774 1217 13299 1232
rect -1774 1211 -1445 1217
rect -1774 255 -1767 1211
rect -1456 255 -1445 1211
rect 13971 1217 15098 1538
rect 15425 1219 15436 1541
rect 15758 1219 15763 1541
rect 15425 1217 15763 1219
rect 15434 1197 15763 1217
rect -1774 226 -1445 255
rect -1774 -623 -1772 226
rect -1449 -623 -1445 226
rect -1774 -654 -1445 -623
rect -1224 982 1544 984
rect -1224 814 14512 982
rect -1224 664 12407 814
rect 13092 664 14512 814
rect -1224 660 14512 664
rect 14852 660 14878 982
rect -1224 655 14878 660
rect -3013 -665 -1441 -654
rect -3013 -1336 -2255 -665
rect -1835 -670 -1441 -665
rect -1835 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -1835 -1336 -1441 -1331
rect -3013 -1341 -1441 -1336
rect -1774 -15992 -1445 -1341
rect -1224 -1544 -895 655
rect 466 653 14878 655
rect 15434 868 15441 1197
rect 14884 618 15213 645
rect -667 444 1547 454
rect -667 125 14656 444
rect -1224 -2224 -1047 -1544
rect -1224 -15428 -895 -2224
rect -667 -14001 -338 125
rect 108 115 14656 125
rect -115 -101 2593 -94
rect -115 -423 14094 -101
rect -115 -13100 214 -423
rect 2416 -430 14094 -423
rect 13765 -1532 14094 -430
rect 13932 -2213 14094 -1532
rect 8399 -7628 8405 -7622
rect 8398 -7698 8405 -7694
rect -115 -13787 42 -13100
rect 200 -13787 214 -13100
rect -667 -14674 -482 -14001
rect -115 -14334 214 -13787
rect 13765 -13979 14094 -2213
rect 14327 -636 14656 115
rect 14499 -1321 14656 -636
rect 13765 -14333 14094 -14312
rect -115 -14347 13267 -14334
rect -115 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -115 -14663 13267 -14484
rect 13646 -14663 13655 -14334
rect 14327 -14517 14656 -1321
rect 14884 -13082 15213 272
rect 15028 -13769 15213 -13082
rect -667 -14889 -338 -14674
rect 14884 -14709 15213 -13769
rect 14327 -14876 14656 -14850
rect -667 -15043 13336 -14889
rect 14002 -15043 14211 -14889
rect -667 -15218 14211 -15043
rect 14645 -15218 14656 -14876
rect 15212 -15053 15213 -14709
rect 14884 -15063 15213 -15053
rect 15212 -15398 15213 -15063
rect 14884 -15418 15213 -15398
rect -1224 -15609 14338 -15428
rect -1224 -15757 886 -15609
rect 1567 -15757 14338 -15609
rect 14772 -15757 14778 -15428
rect 15212 -15757 15213 -15418
rect 15434 -13972 15763 868
rect 15434 -14674 15436 -13972
rect 15747 -13974 15763 -13972
rect 15747 -14654 15766 -13974
rect 15975 -14654 16673 -13974
rect 15747 -14674 15763 -14654
rect 15434 -14694 15763 -14674
rect 15434 -14766 15766 -14694
rect 15521 -14771 15766 -14766
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -14799 15766 -14771
rect 15644 -15986 15646 -14799
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16081 14470 -15993
rect 662 -16090 15766 -16081
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16210 15766 -16204
rect 662 -16313 14469 -16210
rect -1774 -16315 14469 -16313
rect -1774 -16321 10 -16315
rect -9 -16322 10 -16321
rect 661 -16321 14469 -16315
rect 15753 -16321 15766 -16210
rect 10 -17229 661 -16553
<< m234contact >>
rect -1767 255 -1456 1211
rect 13299 1209 13971 1538
rect 15436 1219 15758 1541
rect 12407 664 13092 814
rect 14512 660 14852 987
rect -1816 -1331 -1462 -670
rect 14875 272 15216 618
rect -1047 -2224 -889 -1544
rect 13764 -2213 13932 -1532
rect 42 -13787 200 -13100
rect -482 -14674 -311 -14001
rect 14327 -1321 14499 -636
rect 13757 -14312 14095 -13979
rect 12441 -14484 13126 -14347
rect 13267 -14668 13646 -14333
rect 14872 -13769 15028 -13082
rect 14327 -14850 14665 -14517
rect 13336 -15043 14002 -14877
rect 14877 -15398 15212 -15063
rect 886 -15760 1567 -15609
rect 14338 -15757 14772 -15422
rect 15436 -14674 15747 -13972
rect 15529 -15986 15644 -14771
rect -7 -16313 662 -15992
rect 14468 -16204 15752 -16090
<< m4contact >>
rect 6460 -7395 6484 -7380
rect 6564 -7395 6588 -7380
rect 6668 -7395 6692 -7380
rect 6772 -7395 6796 -7380
rect 6876 -7395 6900 -7380
rect 6980 -7395 7004 -7380
rect 7084 -7395 7108 -7380
rect 7188 -7395 7212 -7380
rect 8405 -7638 8412 -7622
rect 6069 -8380 6093 -8356
rect 6173 -8380 6197 -8356
rect 6277 -8380 6301 -8356
rect 6381 -8380 6405 -8356
rect 6485 -8380 6509 -8356
rect 6589 -8380 6613 -8356
rect 6693 -8380 6717 -8356
rect 6797 -8380 6821 -8356
rect 7121 -8662 7143 -8645
rect 7555 -8662 7577 -8645
rect 7991 -8662 8013 -8645
rect 8424 -8662 8446 -8645
rect 8859 -8662 8881 -8645
rect 9294 -8662 9316 -8645
rect 9726 -8662 9748 -8645
rect 10159 -8662 10181 -8645
<< metal4 >>
rect 13304 1549 13975 2669
rect 1879 1539 15436 1549
rect 15529 1541 15770 1549
rect -1767 1538 15436 1539
rect -1767 1220 13299 1538
rect -1767 1211 8012 1220
rect -1456 1210 8012 1211
rect -1456 255 -1438 1210
rect 13971 1220 15436 1538
rect 13971 1218 13975 1220
rect 15433 1219 15436 1220
rect 15758 1220 15770 1541
rect 15758 1219 15762 1220
rect -1767 -629 -1438 255
rect -1217 984 2672 989
rect -1217 973 14512 984
rect -1217 823 12407 973
rect 13092 823 14512 973
rect -1217 814 14512 823
rect -1217 664 12407 814
rect 13092 664 14512 814
rect -1217 660 14512 664
rect 14852 660 15213 984
rect -1767 -654 -1441 -629
rect -3013 -670 -1441 -654
rect -3013 -1331 -1816 -670
rect -1462 -1331 -1441 -670
rect -3013 -1341 -1441 -1331
rect -1767 -1356 -1441 -1341
rect -1767 -15992 -1438 -1356
rect -1217 -1544 -888 660
rect 1910 655 15213 660
rect 14884 618 15213 655
rect -1217 -1546 -1047 -1544
rect -1217 -2226 -1215 -1546
rect -1057 -2224 -1047 -1546
rect -889 -2224 -888 -1544
rect -1057 -2226 -888 -2224
rect -1217 -15415 -888 -2226
rect -667 451 2201 454
rect -667 443 14656 451
rect -667 127 7141 443
rect 7262 438 14656 443
rect 7262 127 8378 438
rect -667 125 8378 127
rect -667 -13991 -338 125
rect -322 122 8378 125
rect 8499 122 14656 438
rect -667 -14664 -663 -13991
rect -492 -14001 -338 -13991
rect -115 -94 6919 -87
rect -115 -102 14094 -94
rect -115 -103 8177 -102
rect -115 -416 6943 -103
rect -115 -13096 214 -416
rect 2735 -417 6943 -416
rect 7064 -417 8177 -103
rect 2735 -418 8177 -417
rect 8298 -418 14094 -102
rect 2735 -423 14094 -418
rect 13765 -1530 14094 -423
rect 14327 -636 14656 122
rect 14499 -1321 14510 -636
rect 14327 -1323 14510 -1321
rect 13765 -1532 13945 -1530
rect 13932 -2213 13945 -1532
rect 6421 -7395 6460 -7387
rect 7270 -7383 8109 -7378
rect 7212 -7386 8109 -7383
rect 7212 -7391 7278 -7386
rect 6421 -7550 6429 -7395
rect 6564 -7491 6572 -7395
rect 6673 -7448 6679 -7395
rect 6673 -7454 6707 -7448
rect 6701 -7477 6707 -7454
rect 6772 -7463 6780 -7395
rect 6876 -7450 6884 -7395
rect 6980 -7435 6988 -7395
rect 7085 -7418 7093 -7395
rect 7085 -7426 7869 -7418
rect 6980 -7443 7629 -7435
rect 6876 -7458 7389 -7450
rect 6772 -7471 7149 -7463
rect 6701 -7483 6907 -7477
rect 6564 -7499 6669 -7491
rect 6661 -7516 6669 -7499
rect 6901 -7518 6907 -7483
rect 7141 -7518 7149 -7471
rect 7381 -7528 7389 -7458
rect 7621 -7517 7629 -7443
rect 7861 -7518 7869 -7426
rect 8101 -7517 8109 -7386
rect 8412 -7562 8420 -7490
rect 8405 -7570 8420 -7562
rect 8405 -7614 8413 -7570
rect 8405 -7622 8415 -7614
rect 5980 -8347 5989 -8238
rect 5980 -8356 6093 -8347
rect 6183 -8356 6190 -8241
rect 6354 -8260 6363 -8241
rect 6287 -8269 6363 -8260
rect 6287 -8356 6296 -8269
rect 6416 -8334 6423 -8241
rect 6660 -8292 6669 -8241
rect 6390 -8341 6423 -8334
rect 6496 -8301 6669 -8292
rect 6390 -8356 6397 -8341
rect 6496 -8356 6505 -8301
rect 6720 -8318 6729 -8237
rect 6600 -8327 6729 -8318
rect 6600 -8356 6609 -8327
rect 6901 -8333 6909 -8236
rect 6705 -8341 6909 -8333
rect 6705 -8356 6713 -8341
rect 6961 -8357 6969 -8236
rect 8314 -8263 8323 -7704
rect 6821 -8365 6969 -8357
rect 7124 -8272 8323 -8263
rect 7124 -8624 7133 -8272
rect 8314 -8273 8323 -8272
rect 8745 -7778 8749 -7769
rect 8327 -8273 8336 -7783
rect 8747 -7850 8749 -7841
rect 8340 -8273 8349 -7852
rect 8396 -7922 8410 -7914
rect 8402 -7942 8410 -7922
rect 8747 -7926 8749 -7917
rect 8353 -8273 8362 -7954
rect 8366 -7995 8399 -7986
rect 8746 -7994 8749 -7985
rect 8366 -8273 8375 -7995
rect 8379 -8066 8400 -8057
rect 8379 -8273 8388 -8066
rect 8392 -8273 8401 -8139
rect -115 -13778 -111 -13096
rect 28 -13100 214 -13096
rect 28 -13778 42 -13100
rect -115 -13787 42 -13778
rect 200 -13787 214 -13100
rect -492 -14664 -482 -14001
rect -667 -14674 -482 -14664
rect -115 -14334 214 -13787
rect 13765 -13979 14094 -2213
rect -115 -14347 13267 -14334
rect -115 -14484 12441 -14347
rect 13126 -14484 13267 -14347
rect -115 -14532 13267 -14484
rect -115 -14663 12447 -14532
rect 13132 -14663 13267 -14532
rect 13765 -14334 14094 -14312
rect 13646 -14663 14094 -14334
rect 14327 -14517 14656 -1323
rect 14884 -13082 15213 272
rect 15028 -13761 15035 -13082
rect 15212 -13761 15213 -13082
rect 15028 -13769 15213 -13761
rect -667 -14882 -338 -14674
rect -667 -15043 13336 -14882
rect 14327 -14882 14656 -14850
rect 14002 -15043 14656 -14882
rect -667 -15064 14656 -15043
rect 14884 -15063 15213 -13769
rect -667 -15211 13341 -15064
rect 14007 -15211 14656 -15064
rect 15212 -15398 15213 -15063
rect 14884 -15415 15213 -15398
rect -1217 -15421 15213 -15415
rect -1217 -15598 886 -15421
rect 1567 -15422 15213 -15421
rect 1567 -15598 14338 -15422
rect -1217 -15609 14338 -15598
rect -1217 -15744 886 -15609
rect 1567 -15744 14338 -15609
rect 14772 -15744 15213 -15422
rect 15433 -13972 15762 1219
rect 15433 -14674 15436 -13972
rect 15747 -13974 15762 -13972
rect 15747 -14654 16673 -13974
rect 15747 -14674 15762 -14654
rect 15433 -14694 15762 -14674
rect 15433 -14771 15766 -14694
rect 15433 -15986 15529 -14771
rect 15644 -15986 15766 -14771
rect 15433 -15989 15766 -15986
rect 15433 -15992 15768 -15989
rect -1788 -16313 -7 -15992
rect 662 -15993 15768 -15992
rect 662 -16090 15766 -15993
rect 662 -16204 14468 -16090
rect 15752 -16204 15766 -16090
rect 662 -16313 15766 -16204
rect -1788 -16321 15766 -16313
rect -9 -16322 661 -16321
rect 10 -17229 661 -16322
<< m345contact >>
rect 9626 -5342 9649 -5318
rect 9626 -5776 9649 -5752
rect 9626 -6210 9649 -6186
rect 9626 -6644 9649 -6620
rect 9626 -7078 9649 -7054
rect 5614 -7407 5642 -7383
rect 5614 -7511 5642 -7487
rect 9626 -7512 9649 -7488
rect 5614 -7615 5642 -7591
rect 8496 -7602 8504 -7594
rect 9060 -7602 9068 -7594
rect 7650 -7660 7658 -7654
rect 8891 -7662 8899 -7654
rect 7410 -7672 7418 -7666
rect 8495 -7674 8503 -7668
rect 9059 -7674 9067 -7666
rect 5614 -7719 5642 -7695
rect 5614 -7823 5642 -7799
rect 7599 -7804 7607 -7798
rect 5614 -7927 5642 -7903
rect 5614 -8031 5642 -8007
rect 5614 -8135 5642 -8111
rect 8405 -7710 8412 -7694
rect 8871 -7734 8879 -7726
rect 9069 -7746 9077 -7738
rect 8405 -7783 8412 -7768
rect 8636 -7804 8644 -7798
rect 8871 -7806 8879 -7798
rect 9065 -7818 9073 -7810
rect 8640 -7876 8648 -7870
rect 8869 -7878 8877 -7870
rect 8694 -7888 8702 -7882
rect 9067 -7890 9075 -7882
rect 8655 -7948 8663 -7942
rect 8868 -7950 8876 -7942
rect 9626 -7946 9649 -7922
rect 8691 -7960 8699 -7954
rect 9069 -7962 9077 -7954
rect 8640 -8020 8648 -8014
rect 8869 -8022 8877 -8014
rect 9068 -8034 9076 -8026
rect 8689 -8092 8697 -8086
rect 8877 -8094 8885 -8086
rect 8646 -8104 8654 -8098
rect 9067 -8106 9075 -8098
rect 8663 -8164 8671 -8158
rect 8875 -8166 8883 -8158
rect 9626 -8380 9649 -8356
<< m5contact >>
rect 8749 -7638 8758 -7625
rect 8314 -7704 8323 -7695
rect 5848 -7851 5866 -7839
rect 8749 -7710 8758 -7697
rect 8327 -7783 8336 -7770
rect 8749 -7782 8758 -7769
rect 8340 -7852 8349 -7843
rect 8401 -7852 8410 -7843
rect 8749 -7854 8758 -7841
rect 8749 -7926 8758 -7913
rect 8353 -7954 8362 -7945
rect 8402 -7950 8410 -7942
rect 8749 -7998 8758 -7985
rect 8749 -8070 8758 -8057
rect 8749 -8142 8758 -8129
<< metal5 >>
rect 12407 973 13089 2672
rect 12407 661 13089 823
rect 14325 -1320 14510 -640
rect 14657 -1320 16677 -640
rect -3000 -2224 -1215 -1549
rect -1057 -2224 -893 -1549
rect 13759 -2210 13945 -1533
rect 14102 -2210 16674 -1533
rect 9446 -5341 9626 -5328
rect 9446 -5998 9459 -5341
rect 9123 -6011 9459 -5998
rect 9483 -5776 9626 -5766
rect 9483 -5779 9634 -5776
rect 5627 -7462 5635 -7407
rect 5627 -7470 5720 -7462
rect 5630 -7567 5641 -7511
rect 5630 -7578 5694 -7567
rect 5632 -7630 5640 -7615
rect 5632 -7638 5657 -7630
rect 5627 -7783 5635 -7719
rect 5649 -7757 5657 -7638
rect 5683 -7727 5694 -7578
rect 5712 -7684 5720 -7470
rect 9123 -7625 9136 -6011
rect 9483 -6321 9496 -5779
rect 8758 -7638 9136 -7625
rect 9162 -6334 9496 -6321
rect 9540 -6210 9626 -6198
rect 9540 -6211 9637 -6210
rect 5712 -7692 5812 -7684
rect 5683 -7738 5775 -7727
rect 5649 -7765 5747 -7757
rect 5627 -7791 5723 -7783
rect 5623 -7889 5631 -7823
rect 5623 -7897 5696 -7889
rect 5642 -7923 5670 -7918
rect 5632 -8064 5640 -8031
rect 5665 -8051 5670 -7923
rect 5688 -7942 5696 -7897
rect 5715 -7905 5723 -7791
rect 5739 -7870 5747 -7765
rect 5764 -7841 5775 -7738
rect 5804 -7769 5812 -7692
rect 8323 -7704 8405 -7695
rect 9162 -7697 9175 -6334
rect 9540 -6647 9553 -6211
rect 8758 -7710 9175 -7697
rect 9192 -6660 9553 -6647
rect 9619 -6644 9626 -6622
rect 5804 -7777 5866 -7769
rect 8336 -7783 8405 -7770
rect 9192 -7769 9205 -6660
rect 9619 -6960 9632 -6644
rect 8758 -7782 9205 -7769
rect 9244 -6973 9632 -6960
rect 5764 -7851 5848 -7841
rect 9244 -7841 9257 -6973
rect 9620 -7078 9626 -7055
rect 9620 -7281 9633 -7078
rect 5764 -7852 5849 -7851
rect 8349 -7852 8401 -7843
rect 8758 -7854 9257 -7841
rect 9288 -7294 9633 -7281
rect 5739 -7878 5866 -7870
rect 5715 -7913 5866 -7905
rect 9288 -7913 9301 -7294
rect 9618 -7512 9626 -7489
rect 9618 -7602 9631 -7512
rect 8758 -7926 9301 -7913
rect 9322 -7615 9631 -7602
rect 5688 -7950 5866 -7942
rect 8362 -7950 8402 -7942
rect 8362 -7954 8371 -7950
rect 9322 -7985 9335 -7615
rect 9622 -7946 9626 -7932
rect 9622 -7952 9635 -7946
rect 8758 -7998 9335 -7985
rect 9363 -7965 9635 -7952
rect 5665 -8056 5865 -8051
rect 9363 -8057 9376 -7965
rect 5632 -8072 5865 -8064
rect 8758 -8070 9376 -8057
rect 5666 -8113 5866 -8100
rect 5642 -8126 5679 -8113
rect 8758 -8142 9376 -8129
rect 9363 -8350 9376 -8142
rect 9363 -8356 9641 -8350
rect 9363 -8363 9626 -8356
rect -3003 -13778 -111 -13096
rect 28 -13778 209 -13096
rect 14870 -13761 15035 -13086
rect 15212 -13761 16670 -13086
rect 14870 -13764 16670 -13761
rect -3003 -13787 209 -13778
rect -3009 -14664 -663 -13998
rect -492 -14664 -323 -13998
rect -3009 -14672 -323 -14664
rect 12444 -14532 13130 -14343
rect 12444 -14669 12447 -14532
rect 886 -15421 1565 -15415
rect 886 -17232 1565 -15598
rect 12444 -17227 13130 -14669
rect 13339 -15064 14003 -14871
rect 13339 -15230 13341 -15064
rect 13339 -17237 14003 -15230
<< m456contact >>
rect 12407 823 13092 973
rect 7141 127 7262 443
rect 8378 122 8499 438
rect 6943 -417 7064 -103
rect 8177 -418 8298 -102
rect 14510 -1323 14657 -636
rect -1215 -2226 -1057 -1546
rect 13945 -2213 14102 -1530
rect -111 -13778 28 -13096
rect 15035 -13761 15212 -13082
rect -663 -14664 -492 -13991
rect 12447 -14669 13132 -14532
rect 886 -15598 1567 -15421
rect 13341 -15230 14007 -15064
<< m6contact >>
rect 8504 -7602 8512 -7594
rect 9052 -7602 9060 -7594
rect 7658 -7662 7666 -7654
rect 8883 -7662 8891 -7654
rect 7418 -7674 7426 -7666
rect 8503 -7676 8511 -7668
rect 9051 -7674 9059 -7666
rect 8863 -7734 8871 -7726
rect 9061 -7746 9069 -7738
rect 7607 -7806 7615 -7798
rect 8644 -7806 8652 -7798
rect 8863 -7806 8871 -7798
rect 9057 -7818 9065 -7810
rect 8648 -7878 8656 -7870
rect 8861 -7878 8869 -7870
rect 8702 -7890 8710 -7882
rect 9059 -7890 9067 -7882
rect 8663 -7950 8671 -7942
rect 8860 -7950 8868 -7942
rect 8699 -7962 8707 -7954
rect 9061 -7962 9069 -7954
rect 8648 -8022 8656 -8014
rect 8861 -8022 8869 -8014
rect 9060 -8034 9068 -8026
rect 8697 -8094 8705 -8086
rect 8869 -8094 8877 -8086
rect 8654 -8106 8662 -8098
rect 9059 -8106 9067 -8098
rect 8671 -8166 8679 -8158
rect 8867 -8166 8875 -8158
<< metal6 >>
rect 12407 973 13089 2672
rect 12407 661 13089 823
rect 6942 -103 7061 -101
rect 6942 -417 6943 -103
rect -3000 -2224 -1215 -1549
rect -1057 -2224 -893 -1549
rect -3003 -13778 -111 -13096
rect 28 -13778 209 -13096
rect -3003 -13787 209 -13778
rect 6942 -13839 7061 -417
rect 7143 -7666 7262 127
rect 8378 438 8498 442
rect 8178 -102 8298 -101
rect 8178 -7654 8298 -418
rect 7666 -7662 8298 -7654
rect 7143 -7674 7418 -7666
rect 7143 -13829 7262 -7674
rect 8178 -13964 8298 -7662
rect 8378 -13964 8498 122
rect 8841 -7654 8961 -683
rect 8841 -7662 8883 -7654
rect 8891 -7662 8961 -7654
rect 8841 -7726 8961 -7662
rect 8841 -7734 8863 -7726
rect 8871 -7734 8961 -7726
rect 8841 -7798 8961 -7734
rect 8841 -7806 8863 -7798
rect 8871 -7806 8961 -7798
rect 8841 -7870 8961 -7806
rect 8841 -7878 8861 -7870
rect 8869 -7878 8961 -7870
rect 8841 -7942 8961 -7878
rect 8841 -7950 8860 -7942
rect 8868 -7950 8961 -7942
rect 8841 -8014 8961 -7950
rect 8841 -8022 8861 -8014
rect 8869 -8022 8961 -8014
rect 8841 -8086 8961 -8022
rect 8841 -8094 8869 -8086
rect 8877 -8094 8961 -8086
rect 8841 -8158 8961 -8094
rect 8841 -8166 8867 -8158
rect 8875 -8166 8961 -8158
rect -3009 -14664 -663 -13998
rect -492 -14664 -323 -13998
rect 8841 -14229 8961 -8166
rect 9041 -7594 9161 -143
rect 14325 -1320 14510 -640
rect 14657 -1320 16677 -640
rect 13759 -2210 13945 -1533
rect 14102 -2210 16674 -1533
rect 9041 -7602 9052 -7594
rect 9060 -7602 9161 -7594
rect 9041 -7666 9161 -7602
rect 9041 -7674 9051 -7666
rect 9059 -7674 9161 -7666
rect 9041 -7738 9161 -7674
rect 9041 -7746 9061 -7738
rect 9069 -7746 9161 -7738
rect 9041 -7810 9161 -7746
rect 9041 -7818 9057 -7810
rect 9065 -7818 9161 -7810
rect 9041 -7882 9161 -7818
rect 9041 -7890 9059 -7882
rect 9067 -7890 9161 -7882
rect 9041 -7954 9161 -7890
rect 9041 -7962 9061 -7954
rect 9069 -7962 9161 -7954
rect 9041 -8026 9161 -7962
rect 9041 -8034 9060 -8026
rect 9068 -8034 9161 -8026
rect 9041 -8098 9161 -8034
rect 9041 -8106 9059 -8098
rect 9067 -8106 9161 -8098
rect 9041 -14229 9161 -8106
rect 14870 -13761 15035 -13086
rect 15212 -13761 16670 -13086
rect 14870 -13764 16670 -13761
rect -3009 -14672 -323 -14664
rect 12444 -14532 13130 -14343
rect 12444 -14669 12447 -14532
rect 886 -15421 1565 -15415
rect 886 -17232 1565 -15598
rect 12444 -17227 13130 -14669
rect 13339 -15064 14003 -14871
rect 13339 -15230 13341 -15064
rect 13339 -17237 14003 -15230
use pad  pad_48
timestamp 1575998002
transform 1 0 -29 0 1 2000
box -3 -4 672 668
use pad  pad_49
timestamp 1575998002
transform 1 0 860 0 1 2000
box -3 -4 672 668
use pad  pad_50
timestamp 1575998002
transform 1 0 1749 0 1 2000
box -3 -4 672 668
use pad  pad_51
timestamp 1575998002
transform 1 0 2638 0 1 2000
box -3 -4 672 668
use pad  pad_52
timestamp 1575998002
transform 1 0 3527 0 1 2000
box -3 -4 672 668
use pad  pad_53
timestamp 1575998002
transform 1 0 4416 0 1 2000
box -3 -4 672 668
use pad  pad_54
timestamp 1575998002
transform 1 0 5305 0 1 2000
box -3 -4 672 668
use pad  pad_55
timestamp 1575998002
transform 1 0 6194 0 1 2000
box -3 -4 672 668
use pad  pad_56
timestamp 1575998002
transform 1 0 7083 0 1 2000
box -3 -4 672 668
use pad  pad_57
timestamp 1575998002
transform 1 0 7972 0 1 2000
box -3 -4 672 668
use pad  pad_58
timestamp 1575998002
transform 1 0 8861 0 1 2000
box -3 -4 672 668
use pad  pad_59
timestamp 1575998002
transform 1 0 9750 0 1 2000
box -3 -4 672 668
use pad  pad_60
timestamp 1575998002
transform 1 0 10639 0 1 2000
box -3 -4 672 668
use pad  pad_61
timestamp 1575998002
transform 1 0 11528 0 1 2000
box -3 -4 672 668
use pad  pad_62
timestamp 1575998002
transform 1 0 12417 0 1 2000
box -3 -4 672 668
use pad  pad_63
timestamp 1575998002
transform 1 0 13306 0 1 2000
box -3 -4 672 668
use pad  pad_32
timestamp 1575998002
transform 0 1 -2998 -1 0 -662
box -3 -4 672 668
use input_driver  input_driver_0
timestamp 1576123792
transform 0 1 1186 -1 0 -725
box 0 -2 230 102
use pad  pad_16
timestamp 1575998002
transform 0 1 16001 -1 0 -645
box -3 -4 672 668
use pad  pad_33
timestamp 1575998002
transform 0 1 -2998 -1 0 -1551
box -3 -4 672 668
use pad  pad_17
timestamp 1575998002
transform 0 1 16001 -1 0 -1534
box -3 -4 672 668
use pad  pad_34
timestamp 1575998002
transform 0 1 -2998 -1 0 -2440
box -3 -4 672 668
use pad  pad_18
timestamp 1575998002
transform 0 1 16001 -1 0 -2423
box -3 -4 672 668
use pad  pad_35
timestamp 1575998002
transform 0 1 -2998 -1 0 -3329
box -3 -4 672 668
use pad  pad_19
timestamp 1575998002
transform 0 1 16001 -1 0 -3312
box -3 -4 672 668
use pad  pad_36
timestamp 1575998002
transform 0 1 -2998 -1 0 -4218
box -3 -4 672 668
use pad  pad_20
timestamp 1575998002
transform 0 1 16001 -1 0 -4201
box -3 -4 672 668
use pad  pad_37
timestamp 1575998002
transform 0 1 -2998 -1 0 -5107
box -3 -4 672 668
use pad  pad_38
timestamp 1575998002
transform 0 1 -2998 -1 0 -5996
box -3 -4 672 668
use pad  pad_39
timestamp 1575998002
transform 0 1 -2998 -1 0 -6885
box -3 -4 672 668
use pad  pad_40
timestamp 1575998002
transform 0 1 -2998 -1 0 -7774
box -3 -4 672 668
use input_driver  input_driver_3
array 0 0 230 0 7 104
timestamp 1576123792
transform 1 0 5386 0 1 -8169
box 0 -2 230 102
use input_driver  input_driver_2
array 0 0 -230 0 7 104
timestamp 1576123792
transform 0 1 6426 -1 0 -7152
box 0 -2 230 102
use core  core_0
timestamp 1576120818
transform 1 0 6186 0 1 -8168
box -322 -73 2624 656
use input_driver  input_driver_1
array 0 0 230 0 7 -104
timestamp 1576123792
transform 0 -1 6127 1 0 -8608
box 0 -2 230 102
use output_driver  output_driver_0
array 0 0 1098 0 7 434
timestamp 1576124467
transform 1 0 9889 0 1 -8454
box -244 -133 854 301
use pad  pad_21
timestamp 1575998002
transform 0 1 16001 -1 0 -5090
box -3 -4 672 668
use pad  pad_22
timestamp 1575998002
transform 0 1 16001 -1 0 -5979
box -3 -4 672 668
use pad  pad_23
timestamp 1575998002
transform 0 1 16001 -1 0 -6868
box -3 -4 672 668
use pad  pad_24
timestamp 1575998002
transform 0 1 16001 -1 0 -7757
box -3 -4 672 668
use pad  pad_41
timestamp 1575998002
transform 0 1 -2998 -1 0 -8663
box -3 -4 672 668
use pad  pad_42
timestamp 1575998002
transform 0 1 -2998 -1 0 -9552
box -3 -4 672 668
use output_driver  output_driver_1
array 0 0 1098 0 7 434
timestamp 1576124467
transform 0 1 7046 -1 0 -8902
box -244 -133 854 301
use pad  pad_25
timestamp 1575998002
transform 0 1 16001 -1 0 -8646
box -3 -4 672 668
use pad  pad_26
timestamp 1575998002
transform 0 1 16001 -1 0 -9535
box -3 -4 672 668
use pad  pad_43
timestamp 1575998002
transform 0 1 -2998 -1 0 -10441
box -3 -4 672 668
use pad  pad_27
timestamp 1575998002
transform 0 1 16001 -1 0 -10424
box -3 -4 672 668
use pad  pad_44
timestamp 1575998002
transform 0 1 -2998 -1 0 -11330
box -3 -4 672 668
use pad  pad_28
timestamp 1575998002
transform 0 1 16001 -1 0 -11313
box -3 -4 672 668
use pad  pad_45
timestamp 1575998002
transform 0 1 -2998 -1 0 -12219
box -3 -4 672 668
use pad  pad_29
timestamp 1575998002
transform 0 1 16001 -1 0 -12202
box -3 -4 672 668
use pad  pad_46
timestamp 1575998002
transform 0 1 -2998 -1 0 -13108
box -3 -4 672 668
use pad  pad_30
timestamp 1575998002
transform 0 1 16001 -1 0 -13091
box -3 -4 672 668
use pad  pad_47
timestamp 1575998002
transform 0 1 -2998 -1 0 -13997
box -3 -4 672 668
use pad  pad_31
timestamp 1575998002
transform 0 1 16001 -1 0 -13980
box -3 -4 672 668
use pad  pad_0
timestamp 1575998002
transform 1 0 0 0 1 -17223
box -3 -4 672 668
use pad  pad_1
timestamp 1575998002
transform 1 0 889 0 1 -17223
box -3 -4 672 668
use pad  pad_2
timestamp 1575998002
transform 1 0 1778 0 1 -17223
box -3 -4 672 668
use pad  pad_3
timestamp 1575998002
transform 1 0 2667 0 1 -17223
box -3 -4 672 668
use pad  pad_4
timestamp 1575998002
transform 1 0 3556 0 1 -17223
box -3 -4 672 668
use pad  pad_5
timestamp 1575998002
transform 1 0 4445 0 1 -17223
box -3 -4 672 668
use pad  pad_6
timestamp 1575998002
transform 1 0 5334 0 1 -17223
box -3 -4 672 668
use pad  pad_7
timestamp 1575998002
transform 1 0 6223 0 1 -17223
box -3 -4 672 668
use pad  pad_8
timestamp 1575998002
transform 1 0 7112 0 1 -17223
box -3 -4 672 668
use pad  pad_9
timestamp 1575998002
transform 1 0 8001 0 1 -17223
box -3 -4 672 668
use pad  pad_10
timestamp 1575998002
transform 1 0 8890 0 1 -17223
box -3 -4 672 668
use pad  pad_11
timestamp 1575998002
transform 1 0 9779 0 1 -17223
box -3 -4 672 668
use pad  pad_12
timestamp 1575998002
transform 1 0 10668 0 1 -17223
box -3 -4 672 668
use pad  pad_13
timestamp 1575998002
transform 1 0 11557 0 1 -17223
box -3 -4 672 668
use pad  pad_14
timestamp 1575998002
transform 1 0 12446 0 1 -17223
box -3 -4 672 668
use pad  pad_15
timestamp 1575998002
transform 1 0 13335 0 1 -17223
box -3 -4 672 668
<< labels >>
rlabel metal4 6989 -16182 6989 -16182 1 VddIo
rlabel metal4 7131 -15637 7131 -15637 1 GndIo
rlabel metal4 7143 -15058 7143 -15058 1 VddCore
rlabel metal4 7143 -14490 7143 -14490 1 GndCore
<< end >>
