magic
tech scmos
timestamp 1575855885
<< metal1 >>
rect 87 62 91 70
rect 213 62 219 70
rect 207 29 214 40
rect 87 2 92 10
rect 213 2 222 10
<< m3contact >>
rect 164 47 170 53
<< metal3 >>
rect 94 62 207 68
rect 94 42 100 62
rect 144 18 150 21
rect 144 12 213 18
<< metal5 >>
rect 87 51 91 58
use or  or_0
timestamp 1575772227
transform -1 0 133 0 1 -2
box 0 4 42 72
use xor  xor_0
timestamp 1575764352
transform 1 0 121 0 1 -2
box 0 4 62 72
use and  and_0
timestamp 1575855885
transform 1 0 171 0 1 -2
box 0 4 42 72
use mux_4_to_1  mux_4_to_1_0
timestamp 1575855885
transform 1 0 221 0 1 64
box -130 -62 106 6
<< end >>
