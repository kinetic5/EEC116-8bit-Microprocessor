magic
tech scmos
timestamp 1576137657
<< nwell >>
rect -27 131 852 301
rect -20 126 852 131
rect -20 125 39 126
<< pwell >>
rect -20 11 853 12
rect -20 -133 854 11
<< ntransistor >>
rect 47 -80 49 -40
rect 57 -80 59 -40
rect 67 -80 69 -40
rect 77 -80 79 -40
rect 87 -80 89 -40
rect 97 -80 99 -40
rect 107 -80 109 -40
rect 117 -80 119 -40
rect 127 -80 129 -40
rect 137 -80 139 -40
rect 147 -80 149 -40
rect 157 -80 159 -40
rect 167 -80 169 -40
rect 177 -80 179 -40
rect 187 -80 189 -40
rect 197 -80 199 -40
rect 207 -84 209 -38
rect 217 -84 219 -38
rect 227 -84 229 -38
rect 237 -84 239 -38
rect 247 -84 249 -38
rect 257 -84 259 -38
rect 267 -84 269 -38
rect 277 -84 279 -38
rect 287 -84 289 -38
rect 297 -84 299 -38
rect 307 -84 309 -38
rect 317 -84 319 -38
rect 327 -84 329 -38
rect 337 -84 339 -38
rect 347 -84 349 -38
rect 357 -84 359 -38
rect 367 -84 369 -38
rect 377 -84 379 -38
rect 387 -84 389 -38
rect 397 -84 399 -38
rect 407 -84 409 -38
rect 417 -84 419 -38
rect 427 -84 429 -38
rect 437 -84 439 -38
rect 447 -84 449 -38
rect 457 -84 459 -38
rect 467 -84 469 -38
rect 477 -84 479 -38
rect 487 -84 489 -38
rect 497 -84 499 -38
rect 507 -84 509 -38
rect 517 -84 519 -38
rect 527 -84 529 -38
rect 537 -84 539 -38
rect 547 -84 549 -38
rect 557 -84 559 -38
rect 567 -84 569 -38
rect 577 -84 579 -38
rect 587 -84 589 -38
rect 597 -84 599 -38
rect 607 -84 609 -38
rect 617 -84 619 -38
rect 627 -84 629 -38
rect 637 -84 639 -38
rect 647 -84 649 -38
rect 657 -84 659 -38
rect 667 -84 669 -38
rect 677 -84 679 -38
rect 687 -84 689 -38
rect 697 -84 699 -38
rect 707 -84 709 -38
rect 717 -84 719 -38
rect 727 -84 729 -38
rect 737 -84 739 -38
rect 747 -84 749 -38
rect 757 -84 759 -38
rect 767 -84 769 -38
rect 777 -84 779 -38
<< ptransistor >>
rect 47 192 49 252
rect 57 192 59 252
rect 67 192 69 252
rect 77 192 79 252
rect 87 192 89 252
rect 97 192 99 252
rect 107 192 109 252
rect 117 192 119 252
rect 127 192 129 252
rect 137 192 139 252
rect 147 192 149 252
rect 157 192 159 252
rect 167 192 169 252
rect 177 192 179 252
rect 187 192 189 252
rect 197 192 199 252
rect 207 185 209 254
rect 217 185 219 254
rect 227 185 229 254
rect 237 185 239 254
rect 247 185 249 254
rect 257 185 259 254
rect 267 185 269 254
rect 277 185 279 254
rect 287 185 289 254
rect 297 185 299 254
rect 307 185 309 254
rect 317 185 319 254
rect 327 185 329 254
rect 337 185 339 254
rect 347 185 349 254
rect 357 185 359 254
rect 367 185 369 254
rect 377 185 379 254
rect 387 185 389 254
rect 397 185 399 254
rect 407 185 409 254
rect 417 185 419 254
rect 427 185 429 254
rect 437 185 439 254
rect 447 185 449 254
rect 457 185 459 254
rect 467 185 469 254
rect 477 185 479 254
rect 487 185 489 254
rect 497 185 499 254
rect 507 185 509 254
rect 517 185 519 254
rect 527 185 529 254
rect 537 185 539 254
rect 547 185 549 254
rect 557 185 559 254
rect 567 185 569 254
rect 577 185 579 254
rect 587 185 589 254
rect 597 185 599 254
rect 607 185 609 254
rect 617 185 619 254
rect 627 185 629 254
rect 637 185 639 254
rect 647 185 649 254
rect 657 185 659 254
rect 667 185 669 254
rect 677 185 679 254
rect 687 185 689 254
rect 697 185 699 254
rect 707 185 709 254
rect 717 185 719 254
rect 727 185 729 254
rect 737 185 739 254
rect 747 185 749 254
rect 757 185 759 254
rect 767 185 769 254
rect 777 185 779 254
<< ndiffusion >>
rect 46 -80 47 -40
rect 49 -80 50 -40
rect 56 -80 57 -40
rect 59 -80 60 -40
rect 66 -80 67 -40
rect 69 -80 70 -40
rect 76 -80 77 -40
rect 79 -80 80 -40
rect 86 -80 87 -40
rect 89 -80 90 -40
rect 96 -80 97 -40
rect 99 -80 100 -40
rect 106 -80 107 -40
rect 109 -80 110 -40
rect 116 -80 117 -40
rect 119 -80 120 -40
rect 126 -80 127 -40
rect 129 -80 130 -40
rect 136 -80 137 -40
rect 139 -80 140 -40
rect 146 -80 147 -40
rect 149 -80 150 -40
rect 156 -80 157 -40
rect 159 -80 160 -40
rect 166 -80 167 -40
rect 169 -80 170 -40
rect 176 -80 177 -40
rect 179 -80 180 -40
rect 186 -80 187 -40
rect 189 -80 190 -40
rect 196 -80 197 -40
rect 199 -80 200 -40
rect 206 -84 207 -38
rect 209 -84 210 -38
rect 216 -84 217 -38
rect 219 -84 220 -38
rect 226 -84 227 -38
rect 229 -84 230 -38
rect 236 -84 237 -38
rect 239 -84 240 -38
rect 246 -84 247 -38
rect 249 -84 250 -38
rect 256 -84 257 -38
rect 259 -84 260 -38
rect 266 -84 267 -38
rect 269 -84 270 -38
rect 276 -84 277 -38
rect 279 -84 280 -38
rect 286 -84 287 -38
rect 289 -84 290 -38
rect 296 -84 297 -38
rect 299 -84 300 -38
rect 306 -84 307 -38
rect 309 -84 310 -38
rect 316 -84 317 -38
rect 319 -84 320 -38
rect 326 -84 327 -38
rect 329 -84 330 -38
rect 336 -84 337 -38
rect 339 -84 340 -38
rect 346 -84 347 -38
rect 349 -84 350 -38
rect 356 -84 357 -38
rect 359 -84 360 -38
rect 366 -84 367 -38
rect 369 -84 370 -38
rect 376 -84 377 -38
rect 379 -84 380 -38
rect 386 -84 387 -38
rect 389 -84 390 -38
rect 396 -84 397 -38
rect 399 -84 400 -38
rect 406 -84 407 -38
rect 409 -84 410 -38
rect 416 -84 417 -38
rect 419 -84 420 -38
rect 426 -84 427 -38
rect 429 -84 430 -38
rect 436 -84 437 -38
rect 439 -84 440 -38
rect 446 -84 447 -38
rect 449 -84 450 -38
rect 456 -84 457 -38
rect 459 -84 460 -38
rect 466 -84 467 -38
rect 469 -84 470 -38
rect 476 -84 477 -38
rect 479 -84 480 -38
rect 486 -84 487 -38
rect 489 -84 490 -38
rect 496 -84 497 -38
rect 499 -84 500 -38
rect 506 -84 507 -38
rect 509 -84 510 -38
rect 516 -84 517 -38
rect 519 -84 520 -38
rect 526 -84 527 -38
rect 529 -84 530 -38
rect 536 -84 537 -38
rect 539 -84 540 -38
rect 546 -84 547 -38
rect 549 -84 550 -38
rect 556 -84 557 -38
rect 559 -84 560 -38
rect 566 -84 567 -38
rect 569 -84 570 -38
rect 576 -84 577 -38
rect 579 -84 580 -38
rect 586 -84 587 -38
rect 589 -84 590 -38
rect 596 -84 597 -38
rect 599 -84 600 -38
rect 606 -84 607 -38
rect 609 -84 610 -38
rect 616 -84 617 -38
rect 619 -84 620 -38
rect 626 -84 627 -38
rect 629 -84 630 -38
rect 636 -84 637 -38
rect 639 -84 640 -38
rect 646 -84 647 -38
rect 649 -84 650 -38
rect 656 -84 657 -38
rect 659 -84 660 -38
rect 666 -84 667 -38
rect 669 -84 670 -38
rect 676 -84 677 -38
rect 679 -84 680 -38
rect 686 -84 687 -38
rect 689 -84 690 -38
rect 696 -84 697 -38
rect 699 -84 700 -38
rect 706 -84 707 -38
rect 709 -84 710 -38
rect 716 -84 717 -38
rect 719 -84 720 -38
rect 726 -84 727 -38
rect 729 -84 730 -38
rect 736 -84 737 -38
rect 739 -84 740 -38
rect 746 -84 747 -38
rect 749 -84 750 -38
rect 756 -84 757 -38
rect 759 -84 760 -38
rect 766 -84 767 -38
rect 769 -84 770 -38
rect 776 -84 777 -38
rect 779 -84 780 -38
<< pdiffusion >>
rect 46 192 47 252
rect 49 192 50 252
rect 56 192 57 252
rect 59 192 60 252
rect 66 192 67 252
rect 69 192 70 252
rect 76 192 77 252
rect 79 192 80 252
rect 86 192 87 252
rect 89 192 90 252
rect 96 192 97 252
rect 99 192 100 252
rect 106 192 107 252
rect 109 192 110 252
rect 116 192 117 252
rect 119 192 120 252
rect 126 192 127 252
rect 129 192 130 252
rect 136 192 137 252
rect 139 192 140 252
rect 146 192 147 252
rect 149 192 150 252
rect 156 192 157 252
rect 159 192 160 252
rect 166 192 167 252
rect 169 192 170 252
rect 176 192 177 252
rect 179 192 180 252
rect 186 192 187 252
rect 189 192 190 252
rect 196 192 197 252
rect 199 192 200 252
rect 206 185 207 254
rect 209 185 210 254
rect 216 185 217 254
rect 219 185 220 254
rect 226 185 227 254
rect 229 185 230 254
rect 236 185 237 254
rect 239 185 240 254
rect 246 185 247 254
rect 249 185 250 254
rect 256 185 257 254
rect 259 185 260 254
rect 266 185 267 254
rect 269 185 270 254
rect 276 185 277 254
rect 279 185 280 254
rect 286 185 287 254
rect 289 185 290 254
rect 296 185 297 254
rect 299 185 300 254
rect 306 185 307 254
rect 309 185 310 254
rect 316 185 317 254
rect 319 185 320 254
rect 326 185 327 254
rect 329 185 330 254
rect 336 185 337 254
rect 339 185 340 254
rect 346 185 347 254
rect 349 185 350 254
rect 356 185 357 254
rect 359 185 360 254
rect 366 185 367 254
rect 369 185 370 254
rect 376 185 377 254
rect 379 185 380 254
rect 386 185 387 254
rect 389 185 390 254
rect 396 185 397 254
rect 399 185 400 254
rect 406 185 407 254
rect 409 185 410 254
rect 416 185 417 254
rect 419 185 420 254
rect 426 185 427 254
rect 429 185 430 254
rect 436 185 437 254
rect 439 185 440 254
rect 446 185 447 254
rect 449 185 450 254
rect 456 185 457 254
rect 459 185 460 254
rect 466 185 467 254
rect 469 185 470 254
rect 476 185 477 254
rect 479 185 480 254
rect 486 185 487 254
rect 489 185 490 254
rect 496 185 497 254
rect 499 185 500 254
rect 506 185 507 254
rect 509 185 510 254
rect 516 185 517 254
rect 519 185 520 254
rect 526 185 527 254
rect 529 185 530 254
rect 536 185 537 254
rect 539 185 540 254
rect 546 185 547 254
rect 549 185 550 254
rect 556 185 557 254
rect 559 185 560 254
rect 566 185 567 254
rect 569 185 570 254
rect 576 185 577 254
rect 579 185 580 254
rect 586 185 587 254
rect 589 185 590 254
rect 596 185 597 254
rect 599 185 600 254
rect 606 185 607 254
rect 609 185 610 254
rect 616 185 617 254
rect 619 185 620 254
rect 626 185 627 254
rect 629 185 630 254
rect 636 185 637 254
rect 639 185 640 254
rect 646 185 647 254
rect 649 185 650 254
rect 656 185 657 254
rect 659 185 660 254
rect 666 185 667 254
rect 669 185 670 254
rect 676 185 677 254
rect 679 185 680 254
rect 686 185 687 254
rect 689 185 690 254
rect 696 185 697 254
rect 699 185 700 254
rect 706 185 707 254
rect 709 185 710 254
rect 716 185 717 254
rect 719 185 720 254
rect 726 185 727 254
rect 729 185 730 254
rect 736 185 737 254
rect 739 185 740 254
rect 746 185 747 254
rect 749 185 750 254
rect 756 185 757 254
rect 759 185 760 254
rect 766 185 767 254
rect 769 185 770 254
rect 776 185 777 254
rect 779 185 780 254
<< ndcontact >>
rect 40 -80 46 -40
rect 60 -80 66 -40
rect 80 -80 86 -40
rect 100 -80 106 -40
rect 120 -80 126 -40
rect 140 -80 146 -40
rect 160 -80 166 -40
rect 180 -80 186 -40
rect 200 -84 206 -38
rect 220 -84 226 -38
rect 240 -84 246 -38
rect 260 -84 266 -38
rect 280 -84 286 -38
rect 300 -84 306 -38
rect 320 -84 326 -38
rect 340 -84 346 -38
rect 360 -84 366 -38
rect 380 -84 386 -38
rect 400 -84 406 -38
rect 420 -84 426 -38
rect 440 -84 446 -38
rect 460 -84 466 -38
rect 480 -84 486 -38
rect 500 -84 506 -38
rect 520 -84 526 -38
rect 540 -84 546 -38
rect 560 -84 566 -38
rect 580 -84 586 -38
rect 600 -84 606 -38
rect 620 -84 626 -38
rect 640 -84 646 -38
rect 660 -84 666 -38
rect 680 -84 686 -38
rect 700 -84 706 -38
rect 720 -84 726 -38
rect 740 -84 746 -38
rect 760 -84 766 -38
rect 780 -84 786 -38
<< pdcontact >>
rect 40 192 46 252
rect 60 192 66 252
rect 80 192 86 252
rect 100 192 106 252
rect 120 192 126 252
rect 140 192 146 252
rect 160 192 166 252
rect 180 192 186 252
rect 200 185 206 254
rect 220 185 226 254
rect 240 185 246 254
rect 260 185 266 254
rect 280 185 286 254
rect 300 185 306 254
rect 320 185 326 254
rect 340 185 346 254
rect 360 185 366 254
rect 380 185 386 254
rect 400 185 406 254
rect 420 185 426 254
rect 440 185 446 254
rect 460 185 466 254
rect 480 185 486 254
rect 500 185 506 254
rect 520 185 526 254
rect 540 185 546 254
rect 560 185 566 254
rect 580 185 586 254
rect 600 185 606 254
rect 620 185 626 254
rect 640 185 646 254
rect 660 185 666 254
rect 680 185 686 254
rect 700 185 706 254
rect 720 185 726 254
rect 740 185 746 254
rect 760 185 766 254
rect 780 185 786 254
<< psubstratepcontact >>
rect -11 -116 841 -91
<< nsubstratencontact >>
rect -8 263 839 284
<< polysilicon >>
rect 47 252 49 259
rect 57 252 59 259
rect 67 252 69 259
rect 77 252 79 259
rect 87 252 89 259
rect 97 252 99 259
rect 107 252 109 259
rect 117 252 119 259
rect 127 252 129 259
rect 137 252 139 259
rect 147 252 149 259
rect 157 252 159 259
rect 167 252 169 259
rect 177 252 179 259
rect 187 252 189 259
rect 197 252 199 259
rect 207 254 209 259
rect 217 254 219 259
rect 227 254 229 259
rect 237 254 239 259
rect 247 254 249 259
rect 257 254 259 259
rect 267 254 269 259
rect 277 254 279 259
rect 287 254 289 259
rect 297 254 299 259
rect 307 254 309 259
rect 317 254 319 259
rect 327 254 329 259
rect 337 254 339 259
rect 347 254 349 259
rect 357 254 359 259
rect 367 254 369 259
rect 377 254 379 259
rect 387 254 389 259
rect 397 254 399 259
rect 407 254 409 259
rect 417 254 419 259
rect 427 254 429 259
rect 437 254 439 259
rect 447 254 449 259
rect 457 254 459 259
rect 467 254 469 259
rect 477 254 479 259
rect 487 254 489 259
rect 497 254 499 259
rect 507 254 509 259
rect 517 254 519 259
rect 527 254 529 259
rect 537 254 539 259
rect 547 254 549 259
rect 557 254 559 259
rect 567 254 569 259
rect 577 254 579 259
rect 587 254 589 259
rect 597 254 599 259
rect 607 254 609 259
rect 617 254 619 259
rect 627 254 629 259
rect 637 254 639 259
rect 647 254 649 259
rect 657 254 659 259
rect 667 254 669 259
rect 677 254 679 259
rect 687 254 689 259
rect 697 254 699 259
rect 707 254 709 259
rect 717 254 719 259
rect 727 254 729 259
rect 737 254 739 259
rect 747 254 749 259
rect 757 254 759 259
rect 767 254 769 259
rect 777 254 779 259
rect 47 119 49 192
rect 57 119 59 192
rect 67 119 69 192
rect 77 119 79 192
rect 87 119 89 192
rect 97 119 99 192
rect 107 119 109 192
rect 117 119 119 192
rect 127 119 129 192
rect 137 119 139 192
rect 147 119 149 192
rect 157 119 159 192
rect 167 119 169 192
rect 177 119 179 192
rect 187 119 189 192
rect 197 119 199 192
rect 207 119 209 185
rect 217 119 219 185
rect 227 119 229 185
rect 237 119 239 185
rect 247 119 249 185
rect 257 119 259 185
rect 267 119 269 185
rect 277 119 279 185
rect 287 119 289 185
rect 297 119 299 185
rect 307 119 309 185
rect 317 119 319 185
rect 327 119 329 185
rect 337 119 339 185
rect 347 119 349 185
rect 357 119 359 185
rect 367 119 369 185
rect 377 119 379 185
rect 387 119 389 185
rect 397 119 399 185
rect 407 119 409 185
rect 417 119 419 185
rect 427 119 429 185
rect 437 119 439 185
rect 447 119 449 185
rect 457 119 459 185
rect 467 119 469 185
rect 477 119 479 185
rect 487 119 489 185
rect 497 119 499 185
rect 507 119 509 185
rect 517 119 519 185
rect 527 119 529 185
rect 537 119 539 185
rect 547 119 549 185
rect 557 119 559 185
rect 567 119 569 185
rect 577 119 579 185
rect 587 119 589 185
rect 597 119 599 185
rect 607 119 609 185
rect 617 119 619 185
rect 627 119 629 185
rect 637 119 639 185
rect 647 119 649 185
rect 657 119 659 185
rect 667 119 669 185
rect 677 119 679 185
rect 687 119 689 185
rect 697 119 699 185
rect 707 119 709 185
rect 717 119 719 185
rect 727 119 729 185
rect 737 119 739 185
rect 747 119 749 185
rect 757 119 759 185
rect 767 119 769 185
rect 777 119 779 185
rect 787 119 789 259
rect 47 -40 49 30
rect 57 -40 59 30
rect 67 -40 69 30
rect 77 -40 79 30
rect 87 -40 89 30
rect 97 -40 99 30
rect 107 -40 109 30
rect 117 -40 119 30
rect 127 -40 129 30
rect 137 -40 139 30
rect 147 -40 149 30
rect 157 -40 159 30
rect 167 -40 169 30
rect 177 -40 179 30
rect 187 -40 189 30
rect 197 -40 199 30
rect 207 -38 209 30
rect 217 -38 219 30
rect 227 -38 229 30
rect 237 -38 239 30
rect 247 -38 249 30
rect 257 -38 259 30
rect 267 -38 269 30
rect 277 -38 279 30
rect 287 -38 289 30
rect 297 -38 299 30
rect 307 -38 309 30
rect 317 -38 319 30
rect 327 -38 329 30
rect 337 -38 339 30
rect 347 -38 349 30
rect 357 -38 359 30
rect 367 -38 369 30
rect 377 -38 379 30
rect 387 -38 389 30
rect 397 -38 399 30
rect 407 -38 409 30
rect 417 -38 419 30
rect 427 -38 429 30
rect 437 -38 439 30
rect 447 -38 449 30
rect 457 -38 459 30
rect 467 -38 469 30
rect 477 -38 479 30
rect 487 -38 489 30
rect 497 -38 499 30
rect 507 -38 509 30
rect 517 -38 519 30
rect 527 -38 529 30
rect 537 -38 539 30
rect 547 -38 549 30
rect 557 -38 559 30
rect 567 -38 569 30
rect 577 -38 579 30
rect 587 -38 589 30
rect 597 -38 599 30
rect 607 -38 609 30
rect 617 -38 619 30
rect 627 -38 629 30
rect 637 -38 639 30
rect 647 -38 649 30
rect 657 -38 659 30
rect 667 -38 669 30
rect 677 -38 679 30
rect 687 -38 689 30
rect 697 -38 699 30
rect 707 -38 709 30
rect 717 -38 719 30
rect 727 -38 729 30
rect 737 -38 739 30
rect 747 -38 749 30
rect 757 -38 759 30
rect 767 -38 769 30
rect 777 -38 779 30
rect 47 -87 49 -80
rect 57 -87 59 -80
rect 67 -87 69 -80
rect 77 -87 79 -80
rect 87 -87 89 -80
rect 97 -87 99 -80
rect 107 -87 109 -80
rect 117 -87 119 -80
rect 127 -87 129 -80
rect 137 -87 139 -80
rect 147 -87 149 -80
rect 157 -87 159 -80
rect 167 -87 169 -80
rect 177 -87 179 -80
rect 187 -87 189 -80
rect 197 -87 199 -80
rect 207 -87 209 -84
rect 217 -87 219 -84
rect 227 -87 229 -84
rect 237 -87 239 -84
rect 247 -87 249 -84
rect 257 -87 259 -84
rect 267 -87 269 -84
rect 277 -87 279 -84
rect 287 -87 289 -84
rect 297 -87 299 -84
rect 307 -87 309 -84
rect 317 -87 319 -84
rect 327 -87 329 -84
rect 337 -87 339 -84
rect 347 -87 349 -84
rect 357 -87 359 -84
rect 367 -87 369 -84
rect 377 -87 379 -84
rect 387 -87 389 -84
rect 397 -87 399 -84
rect 407 -87 409 -84
rect 417 -87 419 -84
rect 427 -87 429 -84
rect 437 -87 439 -84
rect 447 -87 449 -84
rect 457 -87 459 -84
rect 467 -87 469 -84
rect 477 -87 479 -84
rect 487 -87 489 -84
rect 497 -87 499 -84
rect 507 -87 509 -84
rect 517 -87 519 -84
rect 527 -87 529 -84
rect 537 -87 539 -84
rect 547 -87 549 -84
rect 557 -87 559 -84
rect 567 -87 569 -84
rect 577 -87 579 -84
rect 587 -87 589 -84
rect 597 -87 599 -84
rect 607 -87 609 -84
rect 617 -87 619 -84
rect 627 -87 629 -84
rect 637 -87 639 -84
rect 647 -87 649 -84
rect 657 -87 659 -84
rect 667 -87 669 -84
rect 677 -87 679 -84
rect 687 -87 689 -84
rect 697 -87 699 -84
rect 707 -87 709 -84
rect 717 -87 719 -84
rect 727 -87 729 -84
rect 737 -87 739 -84
rect 747 -87 749 -84
rect 757 -87 759 -84
rect 767 -87 769 -84
rect 777 -87 779 -84
rect 787 -87 789 30
rect 797 -87 799 259
<< polycontact >>
rect 45 30 51 119
rect 55 30 61 119
rect 65 30 71 119
rect 75 30 81 119
rect 85 30 91 119
rect 95 30 101 119
rect 105 30 111 119
rect 115 30 121 119
rect 125 30 131 119
rect 135 30 141 119
rect 145 30 151 119
rect 155 30 161 119
rect 165 30 171 119
rect 175 30 181 119
rect 185 30 191 119
rect 195 30 201 119
rect 215 30 221 119
rect 225 30 231 119
rect 235 30 241 119
rect 245 30 251 119
rect 255 30 261 119
rect 265 30 271 119
rect 275 30 281 119
rect 285 30 291 119
rect 295 30 301 119
rect 305 30 311 119
rect 315 30 321 119
rect 325 30 331 119
rect 335 30 341 119
rect 345 30 351 119
rect 355 30 361 119
rect 365 30 371 119
rect 375 30 381 119
rect 385 30 391 119
rect 395 30 401 119
rect 405 30 411 119
rect 415 30 421 119
rect 425 30 431 119
rect 435 30 441 119
rect 445 30 451 119
rect 455 30 461 119
rect 465 30 471 119
rect 475 30 481 119
rect 485 30 491 119
rect 495 30 501 119
rect 505 30 511 119
rect 515 30 521 119
rect 525 30 531 119
rect 535 30 541 119
rect 545 30 551 119
rect 555 30 561 119
rect 565 30 571 119
rect 575 30 581 119
rect 585 30 591 119
rect 595 30 601 119
rect 605 30 611 119
rect 615 30 621 119
rect 625 30 631 119
rect 635 30 641 119
rect 645 30 651 119
rect 655 30 661 119
rect 665 30 671 119
rect 675 30 681 119
rect 685 30 691 119
rect 695 30 701 119
rect 705 30 711 119
rect 715 30 721 119
rect 725 30 731 119
rect 735 30 741 119
rect 745 30 751 119
rect 755 30 761 119
rect 765 30 771 119
rect 775 30 781 119
rect 785 30 791 119
<< metal1 >>
rect -40 284 841 287
rect -40 263 -8 284
rect 839 263 841 284
rect -40 260 841 263
rect -40 173 31 260
rect 40 252 46 260
rect 60 252 66 260
rect 80 252 86 260
rect 100 252 106 260
rect 120 252 126 260
rect 140 252 146 260
rect 160 252 166 260
rect 180 252 186 260
rect 200 254 206 260
rect 220 254 226 260
rect 240 254 246 260
rect 260 254 266 260
rect 280 254 286 260
rect 300 254 306 260
rect 320 254 326 260
rect 340 254 346 260
rect 360 254 366 260
rect 380 254 386 260
rect 400 254 406 260
rect 420 254 426 260
rect 440 254 446 260
rect 460 254 466 260
rect 480 254 486 260
rect 500 254 506 260
rect 520 254 526 260
rect 540 254 546 260
rect 560 254 566 260
rect 580 254 586 260
rect 600 254 606 260
rect 620 254 626 260
rect 640 254 646 260
rect 660 254 666 260
rect 680 254 686 260
rect 700 254 706 260
rect 720 254 726 260
rect 740 254 746 260
rect 760 254 766 260
rect 780 254 786 260
rect 814 173 841 260
rect -40 142 841 173
rect -40 135 -13 142
rect -16 123 -13 135
rect -16 35 -14 47
rect -41 -2 -14 35
rect 2 30 45 119
rect 51 30 55 119
rect 61 30 65 119
rect 71 30 75 119
rect 81 30 85 119
rect 91 30 95 119
rect 101 30 105 119
rect 111 30 115 119
rect 121 30 125 119
rect 131 30 135 119
rect 141 30 145 119
rect 151 30 155 119
rect 161 30 165 119
rect 171 30 175 119
rect 181 30 185 119
rect 191 30 195 119
rect 201 30 202 119
rect 211 30 215 119
rect 221 30 225 119
rect 231 30 235 119
rect 241 30 245 119
rect 251 30 255 119
rect 261 30 265 119
rect 271 30 275 119
rect 281 30 285 119
rect 291 30 295 119
rect 301 30 305 119
rect 311 30 315 119
rect 321 30 325 119
rect 331 30 335 119
rect 341 30 345 119
rect 351 30 355 119
rect 361 30 365 119
rect 371 30 375 119
rect 381 30 385 119
rect 391 30 395 119
rect 401 30 405 119
rect 411 30 415 119
rect 421 30 425 119
rect 431 30 435 119
rect 441 30 445 119
rect 451 30 455 119
rect 461 30 465 119
rect 471 30 475 119
rect 481 30 485 119
rect 491 30 495 119
rect 501 30 505 119
rect 511 30 515 119
rect 521 30 525 119
rect 531 30 535 119
rect 541 30 545 119
rect 551 30 555 119
rect 561 30 565 119
rect 571 30 575 119
rect 581 30 585 119
rect 591 30 595 119
rect 601 30 605 119
rect 611 30 615 119
rect 621 30 625 119
rect 631 30 635 119
rect 641 30 645 119
rect 651 30 655 119
rect 661 30 665 119
rect 671 30 675 119
rect 681 30 685 119
rect 691 30 695 119
rect 701 30 705 119
rect 711 30 715 119
rect 721 30 725 119
rect 731 30 735 119
rect 741 30 745 119
rect 751 30 755 119
rect 761 30 765 119
rect 771 30 775 119
rect 781 30 785 119
rect -41 -29 841 -2
rect -41 -89 32 -29
rect 40 -89 46 -80
rect 60 -89 66 -80
rect 80 -89 86 -80
rect 100 -89 106 -80
rect 120 -89 126 -80
rect 140 -89 146 -80
rect 160 -89 166 -80
rect 180 -89 186 -80
rect 200 -89 206 -84
rect 220 -89 226 -84
rect 240 -89 246 -84
rect 260 -89 266 -84
rect 280 -89 286 -84
rect 300 -89 306 -84
rect 320 -89 326 -84
rect 340 -89 346 -84
rect 360 -89 366 -84
rect 380 -89 386 -84
rect 400 -89 406 -84
rect 420 -89 426 -84
rect 440 -89 446 -84
rect 460 -89 466 -84
rect 480 -89 486 -84
rect 500 -89 506 -84
rect 520 -89 526 -84
rect 540 -89 546 -84
rect 560 -89 566 -84
rect 580 -89 586 -84
rect 600 -89 606 -84
rect 620 -89 626 -84
rect 640 -89 646 -84
rect 660 -89 666 -84
rect 680 -89 686 -84
rect 700 -89 706 -84
rect 720 -89 726 -84
rect 740 -89 746 -84
rect 760 -89 766 -84
rect 780 -89 786 -84
rect 814 -89 841 -29
rect -41 -91 841 -89
rect -41 -116 -11 -91
<< pm12contact >>
rect 205 30 211 119
<< pdm12contact >>
rect 50 192 56 252
rect 70 192 76 252
rect 90 192 96 252
rect 110 192 116 252
rect 130 192 136 252
rect 150 192 156 252
rect 170 192 176 252
rect 190 192 196 252
rect 210 185 216 254
rect 230 185 236 254
rect 250 185 256 254
rect 270 185 276 254
rect 290 185 296 254
rect 310 185 316 254
rect 330 185 336 254
rect 350 185 356 254
rect 370 185 376 254
rect 390 185 396 254
rect 410 185 416 254
rect 430 185 436 254
rect 450 185 456 254
rect 470 185 476 254
rect 490 185 496 254
rect 510 185 516 254
rect 530 185 536 254
rect 550 185 556 254
rect 570 185 576 254
rect 590 185 596 254
rect 610 185 616 254
rect 630 185 636 254
rect 650 185 656 254
rect 670 185 676 254
rect 690 185 696 254
rect 710 185 716 254
rect 730 185 736 254
rect 750 185 756 254
rect 770 185 776 254
<< ndm12contact >>
rect 50 -80 56 -40
rect 70 -80 76 -40
rect 90 -80 96 -40
rect 110 -80 116 -40
rect 130 -80 136 -40
rect 150 -80 156 -40
rect 170 -80 176 -40
rect 190 -80 196 -40
rect 210 -84 216 -38
rect 230 -84 236 -38
rect 250 -84 256 -38
rect 270 -84 276 -38
rect 290 -84 296 -38
rect 310 -84 316 -38
rect 330 -84 336 -38
rect 350 -84 356 -38
rect 370 -84 376 -38
rect 390 -84 396 -38
rect 410 -84 416 -38
rect 430 -84 436 -38
rect 450 -84 456 -38
rect 470 -84 476 -38
rect 490 -84 496 -38
rect 510 -84 516 -38
rect 530 -84 536 -38
rect 550 -84 556 -38
rect 570 -84 576 -38
rect 590 -84 596 -38
rect 610 -84 616 -38
rect 630 -84 636 -38
rect 650 -84 656 -38
rect 670 -84 676 -38
rect 690 -84 696 -38
rect 710 -84 716 -38
rect 730 -84 736 -38
rect 750 -84 756 -38
rect 770 -84 776 -38
<< metal2 >>
rect 56 192 70 252
rect 76 192 90 252
rect 96 192 110 252
rect 116 192 130 252
rect 136 192 150 252
rect 156 192 170 252
rect 176 192 190 252
rect 196 192 202 252
rect 50 119 202 192
rect 216 185 230 254
rect 236 185 250 254
rect 256 185 270 254
rect 276 185 290 254
rect 296 185 310 254
rect 316 185 330 254
rect 336 185 350 254
rect 356 185 370 254
rect 376 185 390 254
rect 396 185 410 254
rect 416 185 430 254
rect 436 185 450 254
rect 456 185 470 254
rect 476 185 490 254
rect 496 185 510 254
rect 516 185 530 254
rect 536 185 550 254
rect 556 185 570 254
rect 576 185 590 254
rect 596 185 610 254
rect 616 185 630 254
rect 636 185 650 254
rect 656 185 670 254
rect 676 185 690 254
rect 696 185 710 254
rect 716 185 730 254
rect 736 185 750 254
rect 756 185 770 254
rect 776 185 795 254
rect -37 52 -28 118
rect 50 30 205 119
rect 50 -40 202 30
rect 215 -1 795 185
rect 215 -35 813 -1
rect 215 -38 795 -35
rect 56 -80 70 -40
rect 76 -80 90 -40
rect 96 -80 110 -40
rect 116 -80 130 -40
rect 136 -80 150 -40
rect 156 -80 170 -40
rect 176 -80 190 -40
rect 196 -80 202 -40
rect 216 -84 230 -38
rect 236 -84 250 -38
rect 256 -84 270 -38
rect 276 -84 290 -38
rect 296 -84 310 -38
rect 316 -84 330 -38
rect 336 -84 350 -38
rect 356 -84 370 -38
rect 376 -84 390 -38
rect 396 -84 410 -38
rect 416 -84 430 -38
rect 436 -84 450 -38
rect 456 -84 470 -38
rect 476 -84 490 -38
rect 496 -84 510 -38
rect 516 -84 530 -38
rect 536 -84 550 -38
rect 556 -84 570 -38
rect 576 -84 590 -38
rect 596 -84 610 -38
rect 616 -84 630 -38
rect 636 -84 650 -38
rect 656 -84 670 -38
rect 676 -84 690 -38
rect 696 -84 710 -38
rect 716 -84 730 -38
rect 736 -84 750 -38
rect 756 -84 770 -38
rect 776 -84 795 -38
<< m3contact >>
rect 795 -1 840 254
rect 795 -85 813 -35
<< m123contact >>
rect -12 52 2 118
<< metal3 >>
rect -237 84 -234 89
rect -30 52 -12 118
use input_driver  input_driver_0
timestamp 1576130499
transform 1 0 -244 0 1 35
box 0 0 231 100
<< labels >>
rlabel metal1 -31 162 -31 162 1 Vdd
rlabel metal1 -30 7 -30 7 1 Gnd
rlabel m3contact 811 91 811 91 7 out
rlabel metal3 -236 86 -236 86 1 in
<< end >>
