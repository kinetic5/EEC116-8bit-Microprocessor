magic
tech scmos
timestamp 1576128602
<< nwell >>
rect 45 -26 125 11
<< pwell >>
rect 45 -61 125 -26
<< ntransistor >>
rect 69 -38 71 -32
rect 79 -36 81 -32
rect 59 -47 61 -43
rect 99 -40 101 -32
rect 109 -40 111 -32
<< ptransistor >>
rect 59 -9 61 -3
rect 69 -20 71 -14
rect 79 -20 81 -14
rect 99 -20 101 -8
rect 109 -20 111 -8
<< ndiffusion >>
rect 62 -34 69 -32
rect 62 -38 63 -34
rect 68 -38 69 -34
rect 71 -36 73 -32
rect 78 -36 79 -32
rect 81 -36 82 -32
rect 71 -38 75 -36
rect 57 -44 59 -43
rect 52 -47 59 -44
rect 61 -47 67 -43
rect 62 -51 67 -47
rect 98 -40 99 -32
rect 101 -40 102 -32
rect 108 -40 109 -32
rect 111 -40 112 -32
<< pdiffusion >>
rect 62 -3 67 1
rect 58 -9 59 -3
rect 61 -9 67 -3
rect 68 -19 69 -14
rect 62 -20 69 -19
rect 71 -20 73 -14
rect 78 -20 79 -14
rect 81 -20 82 -14
rect 98 -20 99 -8
rect 101 -20 102 -8
rect 108 -20 109 -8
rect 111 -20 112 -8
<< ndcontact >>
rect 52 -44 57 -40
rect 63 -38 68 -34
rect 73 -36 78 -32
rect 92 -40 98 -32
rect 112 -40 118 -32
rect 62 -55 67 -51
<< pdcontact >>
rect 62 1 68 5
rect 52 -9 58 -3
rect 62 -19 68 -14
rect 73 -20 78 -14
rect 92 -20 98 -8
rect 112 -20 118 -8
<< psubstratepcontact >>
rect 49 -58 58 -51
rect 77 -58 86 -51
<< nsubstratencontact >>
rect 49 1 58 7
rect 74 1 85 7
rect 106 1 117 7
<< polysilicon >>
rect 49 -49 51 -1
rect 59 -3 61 0
rect 69 -6 71 -1
rect 79 -5 81 -1
rect 59 -27 61 -9
rect 69 -14 71 -11
rect 79 -14 81 -10
rect 69 -23 71 -20
rect 79 -23 81 -20
rect 59 -43 61 -31
rect 69 -32 71 -29
rect 79 -32 81 -29
rect 69 -41 71 -38
rect 79 -42 81 -36
rect 59 -50 61 -47
rect 69 -49 71 -46
rect 79 -49 81 -47
rect 89 -49 91 -1
rect 99 -8 101 -1
rect 109 -8 111 -1
rect 99 -23 101 -20
rect 109 -23 111 -20
rect 99 -32 101 -29
rect 109 -32 111 -29
rect 99 -49 101 -40
rect 109 -49 111 -40
rect 119 -49 121 -1
<< polycontact >>
rect 57 -31 61 -27
rect 97 -29 103 -23
rect 107 -29 113 -23
<< metal1 >>
rect 45 7 125 9
rect 45 1 49 7
rect 58 5 74 7
rect 58 1 62 5
rect 68 1 74 5
rect 85 1 106 7
rect 117 1 125 7
rect 47 -9 52 -3
rect 58 -9 59 -3
rect 47 -29 53 -9
rect 92 -8 98 1
rect 112 -8 118 1
rect 68 -19 70 -14
rect 52 -34 53 -29
rect 47 -40 53 -34
rect 68 -38 70 -34
rect 73 -23 78 -20
rect 73 -29 97 -23
rect 103 -29 107 -23
rect 73 -32 78 -29
rect 47 -44 52 -40
rect 92 -51 98 -40
rect 112 -51 118 -40
rect 45 -58 49 -51
rect 58 -55 62 -51
rect 67 -55 77 -51
rect 58 -58 77 -55
rect 86 -58 125 -51
rect 45 -59 125 -58
<< pm12contact >>
rect 68 -11 73 -6
rect 77 -10 82 -5
rect 68 -46 73 -41
rect 77 -47 82 -42
<< pdm12contact >>
rect 82 -20 88 -14
rect 102 -20 108 -8
<< ndm12contact >>
rect 82 -38 88 -32
rect 102 -40 108 -32
<< metal2 >>
rect 47 -11 68 -6
rect 47 -29 52 -11
rect 56 -41 61 -27
rect 82 -26 88 -20
rect 82 -32 98 -26
rect 56 -46 68 -41
rect 92 -51 98 -32
<< m3contact >>
rect 82 -10 87 -5
rect 82 -47 87 -42
rect 102 -32 112 -20
<< m123contact >>
rect 47 -34 52 -29
rect 56 -27 61 -22
rect 65 -34 70 -19
<< metal3 >>
rect 56 -10 82 -5
rect 56 -22 61 -10
rect 47 -42 52 -34
rect 47 -47 82 -42
<< labels >>
rlabel nsubstratencontact 109 5 109 5 7 Vdd
rlabel m123contact 58 -25 58 -25 1 enable
rlabel metal2 85 -25 85 -25 1 D
rlabel metal1 75 -27 75 -27 1 mux_out
rlabel metal1 73 -55 73 -55 1 Gnd
<< end >>
