magic
tech scmos
timestamp 1575354951
<< error_p >>
rect 40 51 42 53
<< ntransistor >>
rect 10 28 12 32
rect 30 28 32 32
rect 40 28 42 32
rect 60 28 62 32
<< ptransistor >>
rect 10 44 12 50
rect 30 44 32 50
rect 40 44 42 50
rect 60 44 62 50
<< ndiffusion >>
rect 6 28 10 32
rect 12 28 13 32
rect 29 28 30 32
rect 32 28 40 32
rect 42 28 43 32
rect 59 28 60 32
rect 62 28 66 32
<< pdiffusion >>
rect 6 44 10 50
rect 12 44 16 50
rect 26 48 30 50
rect 29 44 30 48
rect 32 44 40 50
rect 42 48 46 50
rect 42 44 43 48
rect 59 45 60 50
rect 56 44 60 45
rect 62 44 66 50
<< ndcontact >>
rect 13 28 19 32
rect 23 28 29 32
rect 43 28 48 32
<< pdcontact >>
rect 23 44 29 48
rect 43 44 48 48
<< polysilicon >>
rect 0 13 2 55
rect 10 50 12 55
rect 10 43 12 44
rect 10 32 12 38
rect 10 13 12 28
rect 20 13 22 55
rect 30 50 32 51
rect 40 50 42 51
rect 30 41 32 44
rect 40 41 42 44
rect 30 32 32 35
rect 40 32 42 35
rect 30 25 32 28
rect 40 25 42 28
rect 30 13 32 20
rect 40 13 42 21
rect 50 13 52 55
rect 60 50 62 53
rect 60 41 62 44
rect 60 32 62 36
rect 60 13 62 28
rect 70 13 72 55
rect 80 13 82 55
rect 90 13 92 55
rect 100 13 102 55
rect 110 13 112 55
rect 120 13 122 55
<< polycontact >>
rect 40 21 44 25
<< metal1 >>
rect 0 66 122 74
rect 0 2 122 10
<< pm12contact >>
rect 30 51 35 56
rect 10 38 15 43
rect 59 36 64 41
rect 29 20 34 25
<< pdm12contact >>
rect 54 45 59 50
<< ndm12contact >>
rect 54 27 59 32
<< end >>
