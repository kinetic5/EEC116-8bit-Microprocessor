magic
tech scmos
timestamp 1575698634
<< ntransistor >>
rect 10 25 12 29
rect 20 25 22 29
rect 30 25 32 29
rect 50 25 52 29
<< ptransistor >>
rect 10 45 12 51
rect 20 45 22 51
rect 30 45 32 51
rect 50 45 52 51
<< ndiffusion >>
rect 9 25 10 29
rect 12 25 13 29
rect 19 25 20 29
rect 22 25 23 29
rect 29 25 30 29
rect 32 25 33 29
rect 49 25 50 29
rect 52 25 53 29
<< pdiffusion >>
rect 9 45 10 51
rect 12 47 13 51
rect 19 47 20 51
rect 12 45 20 47
rect 22 47 23 51
rect 29 47 30 51
rect 22 45 30 47
rect 32 47 33 51
rect 32 45 39 47
rect 49 45 50 51
rect 52 45 53 51
<< ndcontact >>
rect 3 25 9 29
rect 43 25 49 29
rect 53 25 59 29
<< pdcontact >>
rect 3 45 9 51
rect 43 45 49 51
rect 53 45 59 51
<< polysilicon >>
rect 0 14 2 62
rect 10 51 12 62
rect 20 51 22 62
rect 30 61 32 62
rect 30 51 32 56
rect 10 42 12 45
rect 20 44 22 45
rect 30 40 32 45
rect 10 29 12 33
rect 20 29 22 34
rect 30 29 32 32
rect 10 14 12 25
rect 20 20 22 25
rect 20 14 22 15
rect 30 14 32 25
rect 40 14 42 62
rect 50 51 52 62
rect 50 37 52 45
rect 50 29 52 32
rect 50 14 52 25
rect 60 14 62 62
<< polycontact >>
rect 28 56 34 61
rect 20 38 24 44
rect 28 32 34 36
rect 18 15 24 20
rect 50 32 54 37
<< metal1 >>
rect 0 64 62 72
rect 3 51 9 64
rect 34 56 43 61
rect 53 51 59 64
rect 42 45 43 51
rect 42 44 47 45
rect 24 38 47 44
rect 28 36 34 38
rect 42 29 47 38
rect 3 12 9 25
rect 42 25 43 29
rect 24 15 43 20
rect 53 12 59 25
rect 0 4 62 12
<< m2contact >>
rect 43 55 49 61
rect 50 37 55 42
rect 43 15 49 21
<< pm12contact >>
rect 9 33 14 42
<< pdm12contact >>
rect 13 47 19 53
rect 23 47 29 53
rect 33 47 39 53
<< ndm12contact >>
rect 13 23 19 29
rect 23 23 29 29
rect 33 23 39 29
<< metal2 >>
rect 33 53 39 74
rect 33 42 39 47
rect 14 33 39 42
rect 33 29 39 33
rect 43 61 49 74
rect 43 42 49 55
rect 43 36 50 42
rect 23 2 29 17
rect 43 21 49 36
<< m3contact >>
rect 13 53 19 59
rect 23 53 29 59
rect 13 17 19 23
rect 23 17 29 23
<< metal3 >>
rect 13 23 19 53
rect 23 23 29 53
<< labels >>
rlabel metal1 3 68 3 68 4 Vdd
rlabel metal1 3 8 3 8 2 Gnd
rlabel metal2 36 73 36 73 5 a
rlabel metal2 46 73 46 73 5 b
rlabel metal2 26 3 26 3 1 z
<< end >>
