magic
tech scmos
timestamp 1576013433
<< metal1 >>
rect 1920 494 1931 502
rect 1906 434 1943 442
rect 1918 422 1931 430
rect 1918 362 1930 370
rect 1917 350 1930 358
rect 1917 290 1930 298
rect 1913 278 1930 286
rect 1917 218 1936 226
rect 1914 206 1933 214
rect 1917 146 1930 154
rect 1914 134 1930 142
rect 1910 74 1930 82
rect 1914 62 1930 70
rect 1915 2 1930 10
<< metal2 >>
rect 37 520 43 524
rect -30 514 43 520
rect -213 505 -208 506
rect -13 441 -7 455
rect -13 435 73 441
rect 67 427 73 435
rect 107 431 144 436
rect 139 429 144 431
rect 139 424 148 429
rect -83 389 -74 401
rect 227 369 233 383
rect 227 363 313 369
rect 307 349 313 363
rect 347 359 383 365
rect 377 358 383 359
rect 467 297 473 313
rect 467 291 553 297
rect 547 278 553 291
rect 587 288 624 292
rect 620 279 624 288
rect 707 225 713 239
rect 707 219 793 225
rect 787 206 793 219
rect 827 217 862 221
rect 859 207 863 217
rect 947 153 953 168
rect 947 147 1033 153
rect 1027 133 1033 147
rect 1067 143 1105 148
rect 1100 135 1105 143
rect 1187 69 1193 95
rect 1147 63 1193 69
rect 1236 75 1312 76
rect 1236 74 1309 75
rect 1236 71 1312 74
rect 1236 70 1243 71
rect 1277 70 1312 71
rect 1236 69 1242 70
rect 1247 61 1273 67
rect 1247 44 1253 61
rect 1444 3 1552 9
<< m3contact >>
rect -253 543 -247 549
rect -213 500 -208 505
rect 67 471 73 477
rect 148 424 154 430
rect 307 399 313 405
rect 377 352 383 358
rect -153 317 -145 329
rect 161 317 172 329
rect 547 327 553 333
rect 624 279 630 285
rect 87 245 97 257
rect 403 245 411 257
rect 787 255 793 261
rect 863 207 869 213
rect 1027 183 1033 189
rect 637 176 646 182
rect 1105 135 1111 141
rect 883 101 891 114
rect 1267 111 1273 117
rect 1236 63 1242 69
rect 929 29 937 41
rect 1507 39 1513 45
rect 1439 3 1444 9
<< m123contact >>
rect -180 434 -174 442
<< metal3 >>
rect -243 553 -222 557
rect -95 558 -84 566
rect -287 546 -281 553
rect -243 551 -212 553
rect -247 543 -237 544
rect -297 538 -291 541
rect -253 538 -237 543
rect -228 538 -222 544
rect -218 538 -212 551
rect 12 538 18 552
rect 252 538 258 552
rect 492 538 498 552
rect 732 538 738 552
rect 972 538 978 552
rect 1212 538 1218 552
rect 1452 538 1458 552
rect 1692 538 1698 552
rect 2115 533 2126 545
rect 1950 527 1955 531
rect -180 493 -167 499
rect -180 442 -174 493
rect 225 490 236 494
rect 83 481 98 485
rect 225 486 232 490
rect 33 474 39 481
rect 83 479 108 481
rect 73 471 83 472
rect 23 466 29 469
rect 67 466 83 471
rect 92 464 98 473
rect 102 463 108 479
rect 457 457 467 461
rect 2115 461 2126 473
rect 1950 455 1955 460
rect 154 424 163 430
rect -167 403 -155 410
rect 157 406 163 424
rect 465 419 476 422
rect 323 409 338 413
rect 465 414 477 419
rect 273 402 279 409
rect 323 407 348 409
rect -53 389 -34 401
rect 313 399 329 400
rect 263 394 269 397
rect 307 394 329 399
rect 342 391 348 407
rect 2181 410 2189 627
rect 2193 483 2201 637
rect 2208 555 2216 648
rect 2405 533 2416 545
rect 2240 527 2245 531
rect 2193 472 2216 483
rect 2405 461 2416 473
rect 2240 455 2245 459
rect 2181 402 2205 410
rect 2197 401 2205 402
rect 2115 389 2126 401
rect 1950 383 1955 387
rect 2405 389 2416 401
rect 2240 383 2245 387
rect 383 352 403 358
rect 397 340 403 352
rect 563 337 578 341
rect 705 342 716 350
rect 513 330 519 337
rect 563 335 588 337
rect -145 317 -137 329
rect -123 317 -104 329
rect 172 317 173 329
rect 187 317 206 329
rect 553 327 569 328
rect 503 322 509 324
rect 547 322 569 327
rect -144 302 -137 317
rect 165 311 173 317
rect 582 319 588 335
rect 2115 317 2126 329
rect 1950 311 1955 315
rect 2405 317 2416 329
rect 2240 311 2245 315
rect -144 295 -63 302
rect 690 285 698 290
rect 630 279 643 285
rect -320 247 -313 255
rect -177 240 -174 258
rect -126 246 -95 256
rect 637 261 643 279
rect 803 265 818 269
rect 945 270 956 278
rect 753 258 759 265
rect 803 263 828 265
rect 97 245 102 257
rect 117 245 136 257
rect 96 241 102 245
rect 411 245 413 257
rect 427 245 446 257
rect 793 255 809 256
rect 743 250 749 254
rect 787 250 809 255
rect 407 236 413 245
rect 822 247 828 263
rect 2115 245 2126 257
rect 1950 239 1955 243
rect 2405 245 2416 257
rect 2240 239 2245 243
rect 407 230 410 236
rect 869 207 883 213
rect -176 195 -175 201
rect -167 195 -158 201
rect 455 195 464 206
rect -176 194 -158 195
rect -165 187 -155 194
rect -107 168 -104 186
rect 133 168 136 186
rect 373 168 376 186
rect 877 190 883 207
rect 1043 193 1058 197
rect 1185 198 1196 206
rect 993 186 999 193
rect 1043 191 1068 193
rect 667 173 686 185
rect 1033 183 1049 184
rect 983 178 989 181
rect 1027 178 1049 183
rect 1062 173 1068 191
rect 2115 173 2126 185
rect 1950 167 1955 171
rect 2405 173 2416 185
rect 2240 167 2245 171
rect 1111 135 1123 141
rect 1117 118 1123 135
rect 1283 121 1298 125
rect 1428 126 1436 134
rect 1233 114 1239 121
rect 1283 119 1308 121
rect 891 101 892 114
rect 907 101 926 113
rect 1273 111 1289 112
rect 1223 106 1229 110
rect 1267 106 1289 111
rect 887 92 892 101
rect 1302 101 1308 119
rect 2115 101 2126 113
rect 1950 95 1955 99
rect 2405 101 2416 113
rect 2240 95 2245 99
rect -73 59 72 65
rect -119 43 -115 50
rect -73 41 -67 59
rect -67 32 -63 38
rect -47 30 -34 40
rect 66 24 72 59
rect 297 59 442 65
rect 1177 63 1236 69
rect 1242 63 1244 69
rect 167 39 168 52
rect 297 41 303 59
rect 303 32 307 38
rect 323 30 336 40
rect 436 24 442 59
rect 609 43 625 50
rect 670 24 676 42
rect 1177 45 1183 63
rect 1523 49 1538 53
rect 1668 54 1676 62
rect 1473 42 1479 49
rect 1523 47 1548 49
rect 967 29 986 41
rect 1513 39 1529 40
rect 1463 34 1469 38
rect 1507 34 1529 39
rect 1542 34 1548 47
rect 1897 28 1907 29
rect 2115 29 2126 41
rect 1950 23 1955 27
rect 2405 29 2416 41
rect 2240 23 2245 27
<< m234contact >>
rect 73 533 83 545
rect 313 533 323 545
rect 553 533 563 545
rect 793 533 803 545
rect 1033 533 1043 545
rect 1273 533 1283 545
rect 1513 533 1523 545
rect 1753 533 1763 545
<< m4contact >>
rect -178 568 -170 574
rect -150 568 -142 574
rect -106 568 -99 574
rect -95 566 -84 572
rect -208 545 -202 553
rect -182 536 -173 544
rect -122 536 -113 544
rect -74 543 -64 553
rect -55 535 -48 542
rect -13 533 -3 543
rect 109 546 119 554
rect 139 547 147 554
rect 235 543 243 555
rect 349 546 359 554
rect 379 547 387 554
rect 283 533 293 543
rect 475 543 483 555
rect 589 546 599 554
rect 619 547 627 554
rect 523 533 533 543
rect 715 543 723 555
rect 829 546 839 554
rect 859 547 867 554
rect 763 533 773 543
rect 955 543 963 555
rect 1069 546 1079 554
rect 1099 547 1107 554
rect 1003 533 1013 543
rect 1195 543 1203 555
rect 1309 546 1319 554
rect 1339 547 1347 554
rect 1243 533 1253 543
rect 1435 543 1443 555
rect 1549 546 1559 554
rect 1579 547 1587 554
rect 1483 533 1493 543
rect 1675 543 1683 555
rect 1789 546 1799 554
rect 1819 547 1827 554
rect 1723 533 1733 543
rect 1915 543 1923 555
rect 1937 543 1946 550
rect 2056 547 2065 555
rect -178 506 -170 512
rect -150 506 -142 512
rect -110 506 -102 512
rect 142 496 150 502
rect 179 496 190 502
rect 210 496 221 502
rect -117 463 -108 472
rect -72 463 -63 472
rect 113 475 118 483
rect 137 464 147 472
rect 197 464 207 472
rect 406 471 416 481
rect 425 464 435 474
rect 1937 471 1946 478
rect 2056 475 2065 483
rect 138 434 150 440
rect 210 434 222 440
rect 192 426 198 434
rect 384 424 390 430
rect 422 424 430 430
rect 450 424 458 430
rect -180 403 -167 413
rect -117 402 -109 410
rect 45 390 55 400
rect 123 391 132 400
rect 168 391 177 400
rect 352 403 358 409
rect 378 392 387 400
rect 438 392 447 400
rect 646 399 656 409
rect 665 390 675 400
rect 1937 399 1946 406
rect 2056 403 2065 411
rect 2227 543 2236 550
rect 2498 533 2506 543
rect 2227 471 2236 478
rect 2498 462 2506 472
rect 2227 399 2236 406
rect 2497 390 2505 400
rect 422 360 429 366
rect 622 352 630 357
rect 650 352 658 358
rect 690 352 698 357
rect -234 331 -225 338
rect -187 330 -179 338
rect 123 330 131 338
rect -25 318 -15 328
rect -10 319 -3 327
rect 285 318 295 328
rect 363 319 372 328
rect 410 319 417 328
rect 592 331 598 337
rect 616 320 627 328
rect 677 320 687 328
rect 887 327 896 336
rect 1937 327 1946 334
rect 2056 331 2065 339
rect 905 318 914 327
rect 168 302 176 311
rect 2227 327 2236 334
rect 2207 317 2215 325
rect 2496 318 2504 327
rect -63 295 -56 302
rect 662 285 670 291
rect 862 280 870 286
rect 902 280 910 286
rect 930 280 938 286
rect -234 259 -225 266
rect -136 246 -126 256
rect 53 258 61 266
rect 333 258 343 266
rect 363 258 371 266
rect 215 246 225 256
rect 230 241 243 247
rect 525 246 535 256
rect 603 246 612 255
rect 648 247 657 256
rect 96 229 106 241
rect 832 258 838 264
rect 857 248 867 256
rect 920 248 927 256
rect 1129 255 1136 262
rect 1937 255 1946 262
rect 2056 259 2065 267
rect 1145 245 1155 255
rect 1177 238 1187 245
rect 2227 255 2236 262
rect 2204 246 2212 254
rect 2496 242 2504 251
rect 410 230 418 236
rect 862 217 870 222
rect 901 218 907 224
rect 1102 208 1110 214
rect 1141 208 1150 214
rect 1170 208 1179 214
rect 464 195 474 206
rect 333 186 343 194
rect -250 171 -243 183
rect -25 170 -14 184
rect -10 171 -3 183
rect 212 171 222 182
rect 230 171 237 183
rect 470 183 483 191
rect 573 186 583 194
rect 603 186 611 194
rect 646 176 653 185
rect 765 174 775 184
rect 843 174 852 183
rect 888 175 897 184
rect 1072 186 1078 193
rect 1097 176 1107 184
rect 1157 176 1167 184
rect 1369 183 1376 190
rect 1385 174 1394 184
rect 1937 183 1946 190
rect 2056 187 2065 195
rect 2227 183 2236 190
rect 2205 174 2213 182
rect 2497 175 2505 184
rect 1102 145 1110 150
rect 1142 146 1150 152
rect 1171 146 1179 152
rect 1342 136 1348 142
rect 1378 136 1390 142
rect 714 111 723 120
rect 795 115 805 123
rect 843 114 851 122
rect 1402 126 1408 136
rect 1005 102 1015 112
rect 1083 103 1092 112
rect 1128 103 1137 112
rect 1312 114 1318 121
rect 1336 104 1347 112
rect 1397 104 1407 112
rect 1609 111 1616 118
rect 1625 102 1635 112
rect 1937 111 1946 118
rect 2056 115 2065 123
rect 887 87 897 92
rect 2227 111 2236 118
rect 2206 101 2214 111
rect 2498 101 2506 110
rect -206 39 -197 47
rect 45 26 56 40
rect 1347 66 1353 74
rect 1392 66 1398 74
rect 1402 66 1408 74
rect 1582 64 1590 70
rect 1622 64 1630 70
rect 1650 64 1658 70
rect 143 26 153 40
rect 168 39 177 52
rect 263 42 273 50
rect 410 26 418 40
rect 602 43 609 57
rect 926 56 932 62
rect 515 26 526 40
rect 534 25 543 31
rect 755 26 766 40
rect 771 39 783 47
rect 855 43 865 51
rect 929 41 937 47
rect 1065 30 1075 40
rect 1143 31 1152 40
rect 1188 31 1197 40
rect 1323 31 1332 40
rect 1577 32 1587 40
rect 1637 32 1647 40
rect 1849 39 1856 46
rect 1865 30 1874 40
rect 1937 39 1946 46
rect 2056 43 2065 51
rect 1363 13 1370 21
rect 2227 39 2236 46
rect 2206 29 2214 39
rect 2498 30 2506 39
rect 1529 15 1537 20
rect 1650 2 1658 8
rect 1590 -4 1598 2
rect 1630 -4 1638 2
<< metal4 >>
rect -208 553 -202 578
rect -177 574 -170 588
rect -184 568 -178 574
rect -150 556 -143 568
rect -206 462 -199 496
rect -195 502 -188 553
rect -163 549 -143 556
rect -182 530 -176 536
rect -234 338 -225 351
rect -234 266 -225 279
rect -186 161 -179 330
rect -206 -90 -197 39
rect -188 -11 -181 4
rect -163 -44 -156 549
rect -150 -22 -143 506
rect -136 256 -129 566
rect -117 564 -110 588
rect -106 574 -99 588
rect -90 572 -84 578
rect -117 557 -102 564
rect -120 530 -113 536
rect -109 512 -102 557
rect -94 546 -74 553
rect -110 472 -103 494
rect -108 463 -103 472
rect -116 161 -109 402
rect -117 -33 -110 4
rect -94 3 -87 546
rect -76 543 -74 546
rect -54 530 -48 535
rect -13 528 -3 533
rect -70 472 -63 504
rect -25 328 -18 481
rect 58 400 65 552
rect 76 545 83 649
rect 109 554 115 567
rect 140 554 147 578
rect 235 555 243 584
rect 316 545 323 638
rect 349 554 355 567
rect 380 554 387 578
rect 475 555 483 584
rect 556 545 563 627
rect 589 554 596 567
rect 620 554 627 578
rect 715 555 721 596
rect 796 545 803 616
rect 1036 612 1043 613
rect 829 554 835 567
rect 860 554 867 578
rect 955 555 963 589
rect 1036 545 1043 605
rect 1276 601 1283 613
rect 1069 554 1075 567
rect 1100 554 1107 578
rect 1195 555 1203 584
rect 1276 545 1283 594
rect 1309 554 1315 567
rect 1340 554 1347 578
rect 1435 555 1443 584
rect 1549 554 1555 567
rect 1580 554 1587 578
rect 1675 555 1683 584
rect 1793 554 1799 567
rect 1820 554 1827 578
rect 1915 555 1923 584
rect 2064 578 2065 585
rect 2057 555 2065 578
rect 1931 543 1937 550
rect 142 502 149 505
rect 113 483 117 495
rect 125 400 132 481
rect 137 453 144 464
rect 157 440 164 506
rect 210 502 217 506
rect 150 433 164 440
rect 55 390 65 400
rect -63 278 -56 295
rect -10 298 -3 319
rect -25 161 -14 170
rect -3 -99 4 183
rect 54 161 61 258
rect 97 241 103 292
rect 124 161 131 330
rect 45 -44 56 26
rect 129 26 143 40
rect 129 -22 138 26
rect 145 -11 152 4
rect 157 -33 164 433
rect 170 400 177 466
rect 168 288 174 302
rect 168 -74 177 39
rect 181 -44 188 496
rect 286 475 293 533
rect 197 449 204 464
rect 192 -22 198 426
rect 210 429 218 434
rect 227 388 234 455
rect 384 430 390 460
rect 352 409 358 424
rect 218 256 225 337
rect 288 328 295 409
rect 365 328 372 409
rect 378 382 385 392
rect 230 226 243 241
rect 333 194 341 258
rect 212 -55 222 171
rect 230 -107 237 171
rect 333 142 341 186
rect 364 161 371 258
rect 265 50 273 130
rect 383 -33 390 362
rect 399 3 406 481
rect 428 452 435 464
rect 452 434 458 442
rect 450 430 458 434
rect 410 328 417 392
rect 424 376 430 424
rect 440 387 447 392
rect 440 380 450 387
rect 424 370 438 376
rect 410 236 417 302
rect 410 -33 418 26
rect 422 -22 429 360
rect 433 364 438 370
rect 433 -44 439 364
rect 480 362 486 460
rect 490 400 497 423
rect 526 403 533 533
rect 451 -11 458 356
rect 490 288 496 400
rect 540 301 547 400
rect 552 285 559 434
rect 634 402 646 409
rect 592 337 597 352
rect 620 357 625 358
rect 620 352 622 357
rect 528 256 535 264
rect 605 255 612 337
rect 616 305 623 320
rect 474 198 496 206
rect 463 -33 470 4
rect 474 -104 483 183
rect 488 -66 496 198
rect 573 142 581 186
rect 603 161 610 186
rect 602 57 609 130
rect 515 -11 526 26
rect 534 -68 543 25
rect 612 -11 619 7
rect 623 -33 630 289
rect 634 2 641 402
rect 650 358 658 381
rect 667 380 675 390
rect 698 352 701 357
rect 650 256 657 322
rect 680 305 687 320
rect 694 294 701 352
rect 766 331 773 533
rect 876 329 887 336
rect 646 185 653 229
rect 649 -44 656 7
rect 662 -22 669 285
rect 833 264 837 278
rect 768 184 775 193
rect 845 183 852 265
rect 857 233 864 248
rect 795 123 805 130
rect 843 122 850 154
rect 715 -85 723 111
rect 857 51 865 130
rect 876 113 883 329
rect 907 307 914 318
rect 910 280 916 286
rect 890 184 897 250
rect 877 100 883 113
rect 755 7 766 26
rect 775 -82 783 39
rect 876 2 883 100
rect 887 68 894 87
rect 901 -22 907 218
rect 911 -44 916 280
rect 920 233 927 248
rect 931 231 936 280
rect 931 226 947 231
rect 942 212 947 226
rect 926 62 932 154
rect 929 27 937 41
rect 942 -33 947 207
rect 960 222 966 288
rect 1006 259 1013 533
rect 1115 255 1129 262
rect 960 -11 966 216
rect 1072 193 1077 206
rect 1008 112 1015 120
rect 1085 112 1092 193
rect 1097 164 1104 176
rect 1068 40 1075 49
rect 1093 -11 1099 5
rect 1103 -33 1109 145
rect 1115 2 1122 255
rect 1148 236 1155 245
rect 1154 226 1155 236
rect 1246 187 1253 533
rect 1130 112 1137 176
rect 1159 164 1167 176
rect 1369 151 1376 183
rect 1385 165 1392 174
rect 1142 140 1148 146
rect 1142 134 1162 140
rect 1145 40 1152 121
rect 1143 -44 1149 5
rect 1156 -22 1162 134
rect 1170 -11 1176 146
rect 1374 146 1376 151
rect 1342 142 1348 143
rect 1312 121 1317 134
rect 1190 40 1197 104
rect 1336 92 1343 104
rect 1347 74 1353 94
rect 1323 40 1332 49
rect 1180 -33 1186 5
rect 1335 -11 1341 4
rect 1347 -34 1353 66
rect 1378 50 1384 136
rect 1402 124 1408 126
rect 1388 118 1408 124
rect 1388 102 1393 118
rect 1400 92 1407 104
rect 1378 44 1387 50
rect 1362 13 1363 15
rect 1362 10 1370 13
rect 1381 -45 1387 44
rect 1392 -23 1398 66
rect 1402 -12 1408 66
rect 1412 0 1419 145
rect 1486 115 1493 533
rect 1516 151 1523 533
rect 1505 71 1513 110
rect 1520 69 1525 70
rect 1567 64 1582 70
rect 1520 20 1525 63
rect 1520 15 1529 20
rect 1567 -11 1573 64
rect 1577 16 1584 32
rect 1609 2 1616 111
rect 1626 92 1633 102
rect 1590 -33 1597 -4
rect 1620 64 1622 70
rect 1658 64 1664 70
rect 1620 -44 1626 64
rect 1639 16 1646 32
rect 1657 19 1664 64
rect 1726 43 1733 533
rect 1756 80 1763 533
rect 1931 478 1938 543
rect 2057 483 2065 547
rect 1931 471 1937 478
rect 1911 358 1918 400
rect 1931 406 1938 471
rect 2057 411 2065 475
rect 1931 399 1937 406
rect 1931 334 1938 399
rect 2057 339 2065 403
rect 1931 327 1937 334
rect 1913 296 1920 313
rect 1931 262 1938 327
rect 2057 267 2065 331
rect 1931 255 1937 262
rect 1905 183 1913 242
rect 1931 190 1938 255
rect 2057 195 2065 259
rect 2176 242 2184 593
rect 2189 254 2197 604
rect 2207 325 2215 615
rect 2221 543 2227 550
rect 2221 478 2228 543
rect 2498 514 2506 533
rect 2221 471 2227 478
rect 2221 406 2228 471
rect 2498 444 2506 462
rect 2221 399 2227 406
rect 2221 334 2228 399
rect 2497 400 2505 413
rect 2221 327 2227 334
rect 2221 262 2228 327
rect 2496 327 2504 345
rect 2221 255 2227 262
rect 2189 246 2204 254
rect 2176 234 2205 242
rect 1931 183 1937 190
rect 1931 118 1938 183
rect 2057 123 2065 187
rect 2197 174 2205 234
rect 2221 190 2228 255
rect 2496 251 2504 258
rect 2221 183 2227 190
rect 1931 111 1937 118
rect 1931 46 1938 111
rect 2057 51 2065 115
rect 2206 111 2214 144
rect 2221 118 2228 183
rect 2221 111 2227 118
rect 1657 12 1669 19
rect 1630 -22 1637 -4
rect 1650 -11 1657 2
rect 1662 -33 1669 12
rect 1849 3 1856 39
rect 1867 20 1874 30
rect 1931 39 1937 46
rect 1931 -55 1938 39
rect 2206 39 2214 73
rect 2221 46 2228 111
rect 2221 39 2227 46
rect 2223 30 2236 39
rect 2223 23 2232 30
rect 2223 -65 2236 23
<< m345contact >>
rect -287 553 -278 562
rect -222 553 -213 562
rect -300 529 -291 538
rect -237 536 -228 545
rect -208 496 -199 505
rect -250 391 -243 399
rect -320 319 -313 327
rect -320 241 -307 247
rect -175 195 -167 201
rect -131 43 -119 51
rect 12 552 22 562
rect 43 533 53 543
rect 33 481 42 490
rect -83 453 -76 461
rect -83 389 -74 401
rect 20 457 29 466
rect 2208 648 2216 656
rect 252 552 262 562
rect 2193 637 2201 645
rect 2181 627 2189 634
rect 492 552 502 562
rect 732 552 742 562
rect 972 552 982 562
rect 1212 552 1222 562
rect 1452 552 1462 562
rect 1692 552 1702 562
rect 98 481 107 490
rect 83 464 92 473
rect 93 330 103 338
rect -77 255 -67 266
rect 23 258 32 266
rect 93 186 103 194
rect 225 494 236 500
rect 273 409 282 418
rect 338 409 347 418
rect 260 385 269 394
rect 329 394 338 403
rect 382 362 390 368
rect 457 447 467 457
rect 465 422 476 428
rect 450 356 458 362
rect 513 337 522 346
rect 500 313 509 322
rect 578 337 587 346
rect 569 322 578 331
rect 622 289 630 294
rect 697 379 707 389
rect 705 350 716 356
rect 690 279 698 285
rect 753 265 762 274
rect 818 265 827 274
rect 809 250 818 259
rect 740 241 749 250
rect 937 307 947 317
rect 755 -7 766 7
rect 945 278 956 284
rect 930 216 938 222
rect 993 193 1002 202
rect 1058 193 1067 202
rect 1049 178 1058 187
rect 980 169 989 178
rect 1185 206 1196 212
rect 1417 163 1427 173
rect 1233 121 1242 130
rect 1298 121 1307 130
rect 1289 106 1298 115
rect 1220 97 1229 106
rect 1368 31 1377 40
rect 1428 134 1436 140
rect 1473 49 1482 58
rect 1460 25 1469 34
rect 1538 49 1547 58
rect 1529 34 1538 43
rect 1428 4 1439 9
rect 1657 91 1667 101
rect 1668 62 1676 68
rect 1942 527 1950 534
rect 1960 533 1967 545
rect 2108 533 2115 545
rect 1942 455 1950 462
rect 1960 461 1967 473
rect 2108 461 2115 473
rect 1942 383 1950 390
rect 1960 389 1967 401
rect 2108 389 2115 401
rect 1942 311 1950 318
rect 1960 317 1967 329
rect 2108 317 2115 329
rect 1942 239 1950 246
rect 1960 245 1967 257
rect 2108 245 2115 257
rect 2232 527 2240 534
rect 2250 533 2257 545
rect 2398 533 2405 545
rect 2232 455 2240 462
rect 2250 461 2257 473
rect 2398 461 2405 473
rect 2232 383 2240 390
rect 2250 389 2257 401
rect 2398 389 2405 401
rect 2232 311 2240 318
rect 2250 317 2257 329
rect 2398 317 2405 329
rect 1942 167 1950 174
rect 1960 173 1967 185
rect 2108 173 2115 185
rect 2232 239 2240 246
rect 2250 245 2257 257
rect 2398 245 2405 257
rect 1942 95 1950 102
rect 1960 101 1967 113
rect 2108 101 2115 113
rect 2232 167 2240 174
rect 2250 173 2257 185
rect 2398 173 2405 185
rect 1897 20 1907 28
rect 1942 23 1950 30
rect 1960 29 1967 41
rect 2108 29 2115 41
rect 2232 95 2240 102
rect 2250 101 2257 113
rect 2398 101 2405 113
rect 2232 23 2240 30
rect 2250 29 2257 41
rect 2398 29 2405 41
rect 1927 -62 1938 -55
<< m5contact >>
rect 76 649 83 656
rect -177 588 -170 594
rect -208 578 -202 584
rect -117 588 -110 594
rect -197 553 -188 562
rect -136 566 -121 574
rect -182 521 -173 530
rect -184 506 -178 516
rect -195 493 -186 502
rect -206 453 -197 462
rect -234 351 -225 358
rect -234 279 -225 286
rect -243 171 -233 183
rect -186 154 -179 161
rect -188 -18 -181 -11
rect -152 536 -143 545
rect -90 578 -84 584
rect -122 521 -113 530
rect -112 494 -103 502
rect -116 154 -109 161
rect -150 -29 -143 -22
rect 55 552 65 562
rect -41 538 -32 545
rect -54 521 -46 530
rect -13 518 -3 528
rect -72 504 -63 513
rect -41 506 -32 513
rect -27 481 -18 490
rect 316 638 323 645
rect 140 578 147 585
rect 109 567 116 574
rect 556 627 563 634
rect 380 578 387 585
rect 349 567 356 574
rect 796 616 803 623
rect 620 578 627 584
rect 589 567 596 574
rect 2207 615 2215 623
rect 1036 605 1043 612
rect 860 578 867 585
rect 829 567 836 574
rect 2189 604 2197 612
rect 1276 594 1283 601
rect 1100 578 1107 585
rect 1069 567 1076 574
rect 2176 593 2184 601
rect 1340 578 1347 585
rect 1309 567 1316 574
rect 1580 578 1587 585
rect 1549 567 1556 574
rect 1820 578 1827 585
rect 1793 567 1800 574
rect 2057 578 2064 585
rect 157 506 164 513
rect 113 495 119 501
rect 123 481 132 490
rect 137 444 146 453
rect 210 506 217 513
rect 168 466 177 473
rect -10 290 -3 298
rect 97 292 103 298
rect -63 271 -56 278
rect -25 154 -14 161
rect -94 -7 -84 3
rect -117 -40 -110 -33
rect -163 -51 -156 -44
rect 54 154 61 161
rect 124 154 131 161
rect 145 -18 152 -11
rect 129 -29 138 -22
rect 168 282 174 288
rect 157 -40 164 -33
rect 45 -51 56 -44
rect 284 466 293 475
rect 227 455 234 462
rect 197 442 206 449
rect 210 422 218 429
rect 384 460 390 466
rect 352 424 358 430
rect 286 409 295 418
rect 363 409 372 418
rect 227 381 234 388
rect 216 337 225 346
rect 378 372 388 382
rect 230 218 242 226
rect 192 -29 199 -22
rect 181 -51 188 -44
rect 212 -62 222 -55
rect 364 154 371 161
rect 265 130 273 142
rect 333 130 342 142
rect 480 460 486 466
rect 425 442 435 452
rect 410 392 419 401
rect 442 370 450 380
rect 410 302 417 309
rect 399 -7 406 3
rect 383 -40 390 -33
rect 422 -29 429 -22
rect 410 -40 418 -33
rect 478 356 486 362
rect 490 423 497 430
rect 552 434 559 441
rect 524 394 533 403
rect 540 400 547 407
rect 540 294 547 301
rect 490 282 496 288
rect 592 352 599 358
rect 603 337 612 346
rect 552 278 559 285
rect 528 264 538 274
rect 616 298 626 305
rect 451 -18 458 -11
rect 463 -40 470 -33
rect 433 -51 440 -44
rect 603 154 610 161
rect 573 130 583 142
rect 602 130 609 142
rect 515 -18 526 -11
rect 488 -73 496 -66
rect 612 -18 619 -11
rect 665 370 675 380
rect 648 322 657 329
rect 677 298 687 305
rect 764 322 773 331
rect 694 289 701 294
rect 862 286 871 292
rect 646 229 655 237
rect 634 -7 643 2
rect 623 -40 630 -33
rect 833 278 840 284
rect 843 265 852 274
rect 740 229 749 237
rect 768 193 777 202
rect 857 226 867 233
rect 862 212 870 217
rect 843 154 850 161
rect 795 130 805 142
rect 857 130 865 142
rect 662 -29 669 -22
rect 649 -51 656 -44
rect 905 298 914 307
rect 960 288 966 294
rect 888 250 897 257
rect 887 62 894 68
rect 874 -7 883 2
rect 901 -29 907 -22
rect 920 226 927 233
rect 942 207 947 212
rect 926 154 932 161
rect 929 20 938 27
rect 1004 250 1013 259
rect 960 216 966 222
rect 1072 206 1080 212
rect 1083 193 1092 202
rect 1008 120 1018 130
rect 1097 154 1107 164
rect 1068 49 1077 58
rect 960 -18 966 -11
rect 1093 -18 1099 -11
rect 1144 226 1154 236
rect 1177 230 1187 238
rect 1128 176 1137 185
rect 1244 178 1253 187
rect 1157 154 1167 164
rect 1385 155 1396 165
rect 1143 121 1152 130
rect 1115 -7 1124 2
rect 942 -40 948 -33
rect 1103 -40 1109 -33
rect 1368 145 1374 151
rect 1412 145 1419 151
rect 1312 134 1319 141
rect 1188 104 1197 113
rect 1336 82 1343 92
rect 1347 94 1353 100
rect 1323 49 1332 58
rect 1170 -18 1176 -11
rect 1156 -29 1162 -22
rect 1335 -18 1341 -11
rect 1180 -40 1186 -33
rect 1388 95 1393 102
rect 1398 82 1408 92
rect 1362 4 1370 10
rect 1347 -40 1353 -34
rect 911 -51 917 -44
rect 1143 -51 1149 -44
rect 1516 144 1523 151
rect 1484 106 1493 115
rect 1504 110 1513 119
rect 1491 93 1500 102
rect 1504 62 1513 71
rect 1520 63 1528 69
rect 1412 -7 1421 0
rect 1402 -18 1408 -12
rect 1577 10 1586 16
rect 1623 82 1633 92
rect 1567 -18 1574 -11
rect 1392 -29 1398 -23
rect 1607 -7 1616 2
rect 1590 -40 1598 -33
rect 1637 10 1646 16
rect 1911 400 1918 407
rect 1911 351 1918 358
rect 1913 313 1920 320
rect 1913 289 1920 296
rect 1905 242 1913 250
rect 1905 175 1913 183
rect 2498 504 2506 514
rect 2498 434 2506 444
rect 2497 413 2505 423
rect 2496 345 2504 354
rect 2496 258 2504 267
rect 1756 73 1763 80
rect 2205 144 2214 151
rect 2497 184 2505 193
rect 1724 34 1733 43
rect 1650 -18 1658 -11
rect 1630 -29 1638 -22
rect 2206 73 2214 80
rect 1866 10 1875 20
rect 1847 -7 1856 3
rect 1662 -40 1670 -33
rect 1381 -51 1387 -45
rect 1618 -51 1626 -44
rect 2498 110 2506 124
rect 2498 39 2506 52
rect 2223 -73 2235 -65
<< metal5 >>
rect 83 649 2208 656
rect 76 638 316 645
rect 323 638 2193 645
rect 76 627 556 634
rect 563 627 2181 634
rect 76 616 796 623
rect 803 616 2207 623
rect -162 600 -64 608
rect 76 605 1036 612
rect 1043 605 2189 612
rect -162 598 -110 600
rect -170 588 -117 594
rect -76 590 -64 600
rect 76 594 1276 601
rect 1283 594 2176 601
rect -202 578 -90 584
rect -76 578 109 590
rect 123 585 2064 590
rect 123 578 140 585
rect 147 578 380 585
rect 387 584 860 585
rect 387 578 620 584
rect 627 578 860 584
rect 867 578 1100 585
rect 1107 578 1340 585
rect 1347 578 1580 585
rect 1587 578 1820 585
rect 1827 578 2057 585
rect -121 567 109 574
rect 116 567 349 574
rect 356 567 589 574
rect 596 567 829 574
rect 836 567 1069 574
rect 1076 567 1309 574
rect 1316 567 1549 574
rect 1556 567 1793 574
rect -320 555 -287 562
rect -278 555 -222 562
rect -213 555 -197 562
rect -188 555 12 562
rect 22 555 55 562
rect 65 555 252 562
rect 262 555 492 562
rect 502 555 732 562
rect 742 555 972 562
rect 982 555 1212 562
rect 1222 555 1452 562
rect 1462 555 1692 562
rect 1702 555 1913 562
rect -320 538 -237 545
rect -228 538 -152 545
rect -143 538 -41 545
rect -32 543 53 545
rect -32 538 43 543
rect -173 521 -122 527
rect -113 521 -54 527
rect -178 509 -125 516
rect -41 513 -34 538
rect 1967 533 2108 540
rect 1942 525 1950 527
rect 2257 533 2398 540
rect 2232 525 2240 527
rect -3 518 2410 525
rect -63 506 -41 513
rect 164 507 210 513
rect 1927 504 2498 511
rect 2506 504 2510 511
rect -186 494 -112 501
rect 119 495 225 500
rect -180 483 -27 490
rect -18 483 33 490
rect 42 483 98 490
rect 107 483 123 490
rect 132 483 1920 490
rect -180 466 83 473
rect -197 453 -83 460
rect 92 466 168 473
rect 177 466 284 473
rect 298 472 497 479
rect 298 462 305 472
rect 447 466 471 467
rect 234 455 305 462
rect 390 461 480 466
rect 390 460 453 461
rect 471 460 480 461
rect 490 464 497 472
rect 1927 464 1934 504
rect 490 457 1934 464
rect 146 444 197 449
rect 137 442 197 444
rect 206 442 425 449
rect 1967 461 2108 468
rect 1942 453 1950 455
rect 2257 461 2398 468
rect 2232 453 2240 455
rect 467 447 2410 453
rect 457 446 2410 447
rect 559 434 2498 441
rect 2506 434 2510 441
rect 149 422 210 429
rect 358 428 476 430
rect 358 424 465 428
rect 497 423 2510 430
rect 60 411 273 418
rect 282 411 286 418
rect 295 411 338 418
rect 348 411 363 418
rect 372 411 1913 418
rect -320 391 -250 399
rect 60 394 329 401
rect 338 394 410 401
rect -83 387 -74 389
rect 214 387 227 388
rect -83 381 227 387
rect 419 394 524 401
rect 547 400 1911 407
rect -83 380 221 381
rect 388 372 442 377
rect 394 370 442 372
rect 450 370 665 377
rect 1967 389 2108 396
rect 1942 381 1950 383
rect 2257 389 2398 396
rect 2232 381 2240 383
rect 707 379 2410 381
rect 697 374 2410 379
rect 592 362 716 366
rect -225 351 -179 358
rect 458 356 478 362
rect 592 361 601 362
rect 624 361 716 362
rect 592 358 599 361
rect 705 356 716 361
rect 1918 354 2510 358
rect 1918 351 2496 354
rect 103 330 113 338
rect 225 339 513 346
rect 522 339 578 346
rect 587 339 603 346
rect 612 339 1913 346
rect 2504 351 2510 354
rect 300 322 569 329
rect 578 322 648 329
rect 657 322 764 329
rect 893 321 999 328
rect 893 317 900 321
rect 992 320 999 321
rect 514 310 900 317
rect 514 309 521 310
rect 417 302 521 309
rect 992 313 1913 320
rect 1967 317 2108 324
rect 1942 309 1950 311
rect 2257 317 2398 324
rect 2232 309 2240 311
rect 947 307 2410 309
rect -320 290 -10 298
rect 103 294 540 298
rect 626 298 677 305
rect 687 298 905 305
rect 937 302 2410 307
rect 103 292 547 294
rect 630 289 694 294
rect 862 292 960 294
rect -225 279 -179 286
rect 174 282 490 288
rect 871 288 960 292
rect 1920 289 1944 296
rect 500 278 552 285
rect 618 279 690 284
rect 618 278 698 279
rect 840 278 945 282
rect -56 271 507 278
rect 1937 274 1944 289
rect -320 255 -77 263
rect 32 258 113 266
rect 538 267 753 274
rect 762 267 818 274
rect 828 267 843 274
rect 852 267 1913 274
rect 1937 267 2510 274
rect 540 250 809 257
rect 818 250 888 257
rect 897 250 1004 257
rect 1020 255 1930 263
rect 1132 245 1905 250
rect 756 242 1905 245
rect 1913 242 1930 250
rect 756 237 1140 242
rect 1967 245 2108 252
rect 655 229 740 237
rect 749 229 764 237
rect 867 226 920 233
rect 927 226 1144 233
rect 1942 237 1950 239
rect 2257 245 2398 252
rect 2232 237 2240 239
rect 1187 230 2410 237
rect -320 218 230 226
rect 938 216 960 222
rect 862 207 942 212
rect 1080 206 1185 210
rect -175 194 -167 195
rect 103 186 113 194
rect 777 195 993 202
rect 1002 195 1058 202
rect 1068 195 1083 202
rect 1092 195 1913 202
rect 1926 193 2510 201
rect -320 171 -243 183
rect 780 178 1049 185
rect 1058 178 1128 185
rect 1137 178 1244 185
rect 1926 183 1934 193
rect 1913 175 1934 183
rect -179 154 -116 161
rect -109 154 -25 161
rect -14 154 54 161
rect 61 154 124 161
rect 131 154 364 161
rect 371 154 603 161
rect 610 154 843 161
rect 850 154 926 161
rect 1107 154 1157 161
rect 1167 155 1385 162
rect 1967 173 2108 180
rect 1942 165 1950 167
rect 2257 173 2398 180
rect 2232 165 2240 167
rect 1427 163 2410 165
rect 1417 158 2410 163
rect 1374 145 1412 151
rect 1523 144 2205 151
rect 128 130 265 142
rect 273 130 333 142
rect 342 130 573 142
rect 583 130 602 142
rect 609 130 795 142
rect 805 130 857 142
rect 1319 134 1428 139
rect 1018 123 1143 130
rect 1152 123 1233 130
rect 1242 123 1298 130
rect 1308 123 1913 130
rect 1943 124 2510 132
rect 1943 119 1951 124
rect 1020 106 1188 113
rect 1197 106 1289 113
rect 1298 106 1484 113
rect 1513 111 1951 119
rect 1353 95 1388 101
rect 1500 94 1529 102
rect 1343 82 1398 89
rect 1408 82 1623 89
rect 1967 101 2108 108
rect 1942 93 1950 95
rect 2257 101 2398 108
rect 2232 93 2240 95
rect 1667 91 2410 93
rect 1657 86 2410 91
rect 1763 73 2206 80
rect 894 62 1504 68
rect 1668 69 1676 70
rect 1528 68 1676 69
rect 1528 63 1668 68
rect -162 43 -131 51
rect 1077 51 1323 58
rect 1332 51 1473 58
rect 1482 51 1538 58
rect 1547 51 1920 58
rect 1928 52 2510 58
rect 1928 51 2498 52
rect 1260 40 1529 41
rect 1260 34 1368 40
rect 1377 34 1529 40
rect 1538 34 1724 41
rect 1928 39 1935 51
rect 938 21 1456 27
rect 1854 32 1935 39
rect 1854 27 1861 32
rect 1473 21 1861 27
rect 938 20 1861 21
rect 1967 29 2108 36
rect 1942 21 1950 23
rect 2257 29 2398 36
rect 2506 51 2510 52
rect 2232 21 2240 23
rect 1907 20 2410 21
rect 1449 14 1480 20
rect -320 -7 -94 0
rect -84 -7 399 0
rect 406 -7 634 0
rect 643 -7 755 0
rect 1586 10 1637 16
rect 1646 10 1866 16
rect 1897 14 2410 20
rect 1370 4 1428 9
rect 766 -7 874 0
rect 883 -7 1115 0
rect 1124 -7 1412 0
rect 1421 -7 1607 0
rect 1616 -7 1847 0
rect -320 -18 -188 -11
rect -181 -18 145 -11
rect 152 -18 451 -11
rect 458 -18 515 -11
rect 526 -18 612 -11
rect 619 -18 960 -11
rect 966 -18 1093 -11
rect 1099 -18 1170 -11
rect 1176 -18 1335 -11
rect 1341 -12 1567 -11
rect 1341 -18 1402 -12
rect 1408 -18 1567 -12
rect 1574 -18 1650 -11
rect 1658 -18 1920 -11
rect -320 -29 -150 -22
rect -143 -29 129 -22
rect 138 -29 192 -22
rect 199 -29 422 -22
rect 429 -29 662 -22
rect 669 -29 901 -22
rect 907 -29 1156 -22
rect 1162 -23 1630 -22
rect 1162 -29 1392 -23
rect 1398 -29 1630 -23
rect 1638 -29 1920 -22
rect -320 -40 -117 -33
rect -110 -40 157 -33
rect 164 -40 383 -33
rect 390 -40 410 -33
rect 418 -40 463 -33
rect 470 -40 623 -33
rect 630 -40 942 -33
rect 948 -40 1103 -33
rect 1109 -40 1180 -33
rect 1186 -34 1590 -33
rect 1186 -40 1347 -34
rect 1353 -40 1590 -34
rect 1598 -40 1662 -33
rect 1670 -40 1920 -33
rect -320 -51 -163 -44
rect -156 -51 45 -44
rect 56 -51 181 -44
rect 188 -51 433 -44
rect 440 -51 649 -44
rect 656 -51 911 -44
rect 917 -51 1143 -44
rect 1149 -45 1618 -44
rect 1149 -51 1381 -45
rect 1387 -51 1618 -45
rect 1626 -51 1920 -44
rect 222 -62 1927 -55
rect 496 -73 2223 -66
<< m456contact >>
rect -106 588 -97 596
rect -197 566 -184 574
rect 134 505 149 513
rect 440 434 452 442
rect -179 413 -167 423
rect 646 381 658 390
rect 605 350 620 358
rect 1098 214 1110 222
rect 1141 214 1153 222
rect 1167 214 1179 222
rect 1336 143 1348 151
rect -191 4 -181 13
rect -117 4 -107 13
rect 142 4 152 13
rect 462 4 470 12
rect 610 7 619 15
rect 649 7 658 15
rect 1091 5 1099 13
rect 1141 5 1149 13
rect 1180 5 1188 13
rect 1335 4 1343 12
<< m6contact >>
rect -180 598 -162 608
rect 109 578 123 590
rect -125 506 -114 517
rect 136 422 149 430
rect -179 350 -167 358
rect 113 330 123 338
rect -179 278 -167 286
rect 610 278 618 286
rect 113 258 123 266
rect -179 186 -167 194
rect 113 186 123 194
rect 116 130 128 146
rect -174 43 -162 51
<< metal6 >>
rect -180 591 -167 598
rect -191 13 -184 566
rect -174 423 -167 591
rect -106 513 -99 588
rect -114 506 -99 513
rect -174 358 -167 413
rect -174 286 -167 350
rect -174 194 -167 278
rect -174 51 -167 186
rect -114 13 -107 506
rect 116 338 123 578
rect 142 430 149 505
rect 116 266 123 330
rect 116 194 123 258
rect 116 146 123 186
rect 142 13 149 422
rect 440 12 448 434
rect 610 286 617 350
rect 610 15 617 278
rect 651 15 658 381
rect 930 41 938 325
rect 440 4 462 12
rect 1102 13 1110 214
rect 1099 5 1110 13
rect 1141 13 1149 214
rect 1167 13 1175 214
rect 1167 5 1180 13
rect 1341 12 1348 143
rect 1343 4 1348 12
use logic  logic_0
timestamp 1576013433
transform 1 0 -407 0 1 504
box 85 2 327 70
use two_1_mux  two_1_mux_0
timestamp 1576013433
transform 1 0 -125 0 1 565
box 45 -59 125 9
use fadder  fadder_0
timestamp 1576013433
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1576013433
transform 1 0 -87 0 1 432
box 85 2 327 70
use inputff  inputff_0
timestamp 1576013433
transform 1 0 -174 0 1 482
box -76 -120 134 -52
use driver  driver_0
timestamp 1576013433
transform 1 0 -32 0 1 421
box -8 -59 92 9
use fadder  fadder_1
timestamp 1576013433
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1576013433
transform 1 0 153 0 1 360
box 85 2 327 70
use inputff  inputff_1
timestamp 1576013433
transform 1 0 -244 0 1 410
box -76 -120 134 -52
use driver  driver_1
timestamp 1576013433
transform 1 0 -102 0 1 349
box -8 -59 92 9
use inputff  inputff_2
timestamp 1576013433
transform 1 0 66 0 1 410
box -76 -120 134 -52
use driver  driver_2
timestamp 1576013433
transform 1 0 208 0 1 349
box -8 -59 92 9
use fadder  fadder_2
timestamp 1576013433
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1576013433
transform 1 0 393 0 1 288
box 85 2 327 70
use dff  dff_0
timestamp 1576013433
transform 1 0 -320 0 1 279
box 0 -61 150 7
use driver  driver_8
timestamp 1576013433
transform 1 0 -172 0 1 277
box -8 -59 92 9
use inputff  inputff_3
timestamp 1576013433
transform 1 0 -4 0 1 338
box -76 -120 134 -52
use driver  driver_3
timestamp 1576013433
transform 1 0 138 0 1 277
box -8 -59 92 9
use inputff  inputff_4
timestamp 1576013433
transform 1 0 306 0 1 338
box -76 -120 134 -52
use driver  driver_4
timestamp 1576013433
transform 1 0 448 0 1 277
box -8 -59 92 9
use fadder  fadder_3
timestamp 1576013433
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1576013433
transform 1 0 633 0 1 216
box 85 2 327 70
use dff  dff_3
timestamp 1576013433
transform 1 0 -250 0 1 207
box 0 -61 150 7
use driver  driver_11
timestamp 1576013433
transform 1 0 -102 0 1 205
box -8 -59 92 9
use dff  dff_2
timestamp 1576013433
transform 1 0 -10 0 1 207
box 0 -61 150 7
use driver  driver_10
timestamp 1576013433
transform 1 0 138 0 1 205
box -8 -59 92 9
use dff  dff_1
timestamp 1576013433
transform 1 0 230 0 1 207
box 0 -61 150 7
use driver  driver_9
timestamp 1576013433
transform 1 0 378 0 1 205
box -8 -59 92 9
use inputff  inputff_5
timestamp 1576013433
transform 1 0 546 0 1 266
box -76 -120 134 -52
use driver  driver_5
timestamp 1576013433
transform 1 0 688 0 1 205
box -8 -59 92 9
use fadder  fadder_4
timestamp 1576013433
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1576013433
transform 1 0 873 0 1 144
box 85 2 327 70
use inputff  inputff_6
timestamp 1576013433
transform 1 0 786 0 1 194
box -76 -120 134 -52
use driver  driver_6
timestamp 1576013433
transform 1 0 928 0 1 133
box -8 -59 92 9
use fadder  fadder_5
timestamp 1576013433
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1576013433
transform 1 0 1113 0 1 72
box 85 2 327 70
use dff  dff_6
timestamp 1576013433
transform 1 0 -210 0 1 63
box 0 -61 150 7
use inv_9_6  inv_9_6_2
timestamp 1576013433
transform 1 0 -70 0 1 62
box 0 -60 30 8
use driver  driver_15
timestamp 1576013433
transform 1 0 -32 0 1 61
box -8 -59 92 9
use driver  driver_16
timestamp 1576013433
transform 1 0 68 0 1 61
box -8 -59 92 9
use dff  dff_5
timestamp 1576013433
transform 1 0 160 0 1 63
box 0 -61 150 7
use inv_9_6  inv_9_6_1
timestamp 1576013433
transform 1 0 300 0 1 62
box 0 -60 30 8
use driver  driver_13
timestamp 1576013433
transform 1 0 338 0 1 61
box -8 -59 92 9
use driver  driver_14
timestamp 1576013433
transform 1 0 438 0 1 61
box -8 -59 92 9
use dff  dff_4
timestamp 1576013433
transform 1 0 530 0 1 63
box 0 -61 150 7
use driver  driver_12
timestamp 1576013433
transform 1 0 678 0 1 61
box -8 -59 92 9
use inputff  inputff_7
timestamp 1576013433
transform 1 0 846 0 1 122
box -76 -120 134 -52
use driver  driver_7
timestamp 1576013433
transform 1 0 988 0 1 61
box -8 -59 92 9
use fadder  fadder_6
timestamp 1576013433
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1576013433
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1576013433
transform 1 0 1353 0 1 0
box 85 2 327 70
use enff  enff_0
array 0 0 191 0 7 72
timestamp 1576013433
transform 1 0 1973 0 1 2
box -43 0 147 68
use driver  driver_17
array 0 0 100 0 7 72
timestamp 1576013433
transform 1 0 2128 0 1 61
box -8 -59 92 9
use enff  enff_1
array 0 0 190 0 7 72
timestamp 1576013433
transform 1 0 2263 0 1 2
box -43 0 147 68
use driver  driver_18
array 0 0 100 0 7 72
timestamp 1576013433
transform 1 0 2418 0 1 61
box -8 -59 92 9
use mult  mult_0
timestamp 1576013433
transform 1 0 241 0 1 432
box -241 -432 1689 142
<< labels >>
rlabel m4contact 430 469 430 469 1 4mux_to_2mux_1
rlabel m4contact -8 535 -8 535 1 nz0
rlabel metal5 1659 88 1659 88 1 nz6
rlabel m345contact 459 448 459 448 1 nz1
rlabel m345contact 700 380 700 380 1 nz2
rlabel m345contact 941 308 941 308 1 nz3
rlabel m5contact 1181 233 1181 233 1 nz4
rlabel metal5 1420 160 1420 160 1 nz5
rlabel m5contact 1824 582 1824 582 1 clk
rlabel metal4 239 580 239 580 1 x0
rlabel metal4 1439 580 1439 580 1 x5
rlabel metal4 1679 581 1679 581 1 x6
rlabel metal4 1920 581 1920 581 1 x7
rlabel metal4 1199 581 1199 581 1 x4
rlabel metal4 959 580 959 580 1 x3
rlabel metal4 718 590 718 590 1 x2
rlabel metal4 479 576 479 576 1 x1
rlabel metal3 -318 251 -318 251 3 Actrl
rlabel m5contact -238 177 -238 177 1 Bctrl
rlabel metal4 538 24 538 24 1 opcode2
rlabel metal5 1640 -3 1640 -3 1 _op2
rlabel metal5 1639 -15 1639 -15 1 _op1
rlabel metal5 1639 -26 1639 -26 1 _op0
rlabel metal5 1639 -37 1639 -37 1 _nop1
rlabel metal5 1639 -48 1639 -48 1 _nop0
rlabel m4contact 170 49 170 49 1 opcode1
rlabel metal4 -204 36 -204 36 1 opcode0
rlabel metal4 57 395 57 395 1 _y0
rlabel m345contact -246 395 -246 395 1 y0
rlabel m4contact -20 322 -20 322 1 _y1
rlabel m345contact -317 323 -317 323 3 y1
rlabel m4contact 291 322 291 322 1 _y2
rlabel m4contact -6 323 -6 323 1 y2
rlabel m345contact -72 260 -72 260 1 y3
rlabel m4contact 220 251 220 251 1 _y3
rlabel metal4 238 240 238 240 1 y4
rlabel m5contact 534 270 534 270 1 _y4
rlabel metal4 476 180 476 180 1 y5
rlabel m5contact 773 198 773 198 1 _y5
rlabel metal4 716 109 716 109 1 y6
rlabel m5contact 1013 125 1013 125 1 _y6
rlabel m5contact 1073 54 1073 54 1 _y7
rlabel metal4 776 38 776 38 1 y7
rlabel metal4 -203 489 -203 489 1 _s0
rlabel metal4 1934 546 1934 546 1 c_en
rlabel metal5 1972 321 1972 321 1 z3
rlabel metal5 1972 392 1972 392 1 z2
rlabel metal5 1972 465 1972 465 1 z1
rlabel metal5 1972 537 1972 537 1 z0
rlabel metal5 1972 248 1972 248 1 z4
rlabel metal5 1972 176 1972 176 1 z5
rlabel metal5 1972 105 1972 105 1 z6
rlabel metal5 1900 17 1900 17 1 nz7
rlabel metal5 1918 36 1918 36 1 d7
rlabel metal5 1918 115 1918 115 1 d6
rlabel m5contact 1917 316 1917 316 1 d4
rlabel m5contact 1914 404 1914 404 1 d3
rlabel metal5 1903 437 1903 437 1 d1
rlabel metal5 1916 460 1916 460 1 d0
rlabel metal5 1915 427 1915 427 1 d2
rlabel metal5 2117 652 2117 652 5 c0
rlabel metal5 2117 641 2117 641 1 c1
rlabel metal5 2117 630 2117 630 1 c2
rlabel metal5 2117 619 2117 619 1 c3
rlabel metal5 2117 608 2117 608 1 c4
rlabel metal5 2117 598 2117 598 1 c5
rlabel metal5 1926 246 1926 246 1 d5
rlabel metal4 2224 546 2224 546 1 d_en
rlabel m4contact -7 177 -7 177 1 Cen
rlabel metal4 232 169 232 169 1 Den
<< end >>
