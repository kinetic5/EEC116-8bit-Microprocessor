magic
tech scmos
timestamp 1575849300
<< metal3 >>
rect -163 553 -141 557
rect -207 546 -201 553
rect -163 551 -132 553
rect -138 538 -132 551
rect 12 538 18 552
rect 252 538 258 552
rect 492 538 498 552
rect 732 538 738 552
rect 972 538 978 552
rect 1212 538 1218 552
rect 1452 538 1458 552
rect 1692 538 1698 552
rect 83 481 99 485
rect 33 474 39 481
rect 83 479 108 481
rect 102 463 108 479
rect 323 409 339 413
rect 273 402 279 409
rect 323 407 348 409
rect 342 391 348 407
rect 563 337 579 341
rect 513 330 519 337
rect 563 335 588 337
rect 582 319 588 335
rect 803 265 819 269
rect 753 258 759 265
rect 803 263 828 265
rect 822 247 828 263
rect 1043 193 1059 197
rect 993 186 999 193
rect 1043 191 1068 193
rect 1062 173 1068 191
rect 1283 121 1299 125
rect 1233 114 1239 121
rect 1283 119 1308 121
rect 1302 101 1308 119
rect 1523 49 1539 53
rect 1473 42 1479 49
rect 1523 47 1548 49
rect 1542 34 1548 47
<< m4contact >>
rect -117 463 -108 472
rect -72 463 -63 472
rect 123 391 132 400
rect 363 318 372 327
rect 603 246 612 255
rect 843 174 852 183
rect 1083 102 1092 111
rect 1143 31 1152 40
rect 1323 31 1332 40
<< metal4 >>
rect -117 472 -108 553
rect 123 400 132 481
rect 363 327 372 409
rect 603 255 612 337
rect 843 183 852 265
rect 1083 111 1092 193
rect 1143 40 1152 121
rect 1323 40 1332 49
<< m345contact >>
rect -207 553 -198 562
rect -141 553 -132 562
rect 12 552 22 562
rect 252 552 262 562
rect 492 552 502 562
rect 732 552 742 562
rect 972 552 982 562
rect 1212 552 1222 562
rect 1452 552 1462 562
rect 1692 552 1702 562
rect 46 533 56 543
rect 286 533 296 543
rect 526 533 536 543
rect 766 533 776 543
rect 1006 533 1016 543
rect 1246 533 1256 543
rect 1726 533 1736 543
rect 33 481 42 490
rect 99 481 108 490
rect 273 409 282 418
rect 339 409 348 418
rect 513 337 522 346
rect 579 337 588 346
rect 753 265 762 274
rect 819 265 828 274
rect 993 193 1002 202
rect 1059 193 1068 202
rect 1233 121 1242 130
rect 1299 121 1308 130
rect 1473 49 1482 58
rect 1539 49 1548 58
<< m5contact >>
rect -117 553 -108 562
rect 123 481 132 490
rect 363 409 372 418
rect 603 337 612 346
rect 843 265 852 274
rect 1083 193 1092 202
rect 1143 121 1152 130
rect 1323 49 1332 58
<< metal5 >>
rect -180 483 0 490
rect 60 411 240 418
rect 300 339 480 346
rect 540 267 720 274
rect 780 195 960 202
rect 1020 123 1143 130
rect 1152 123 1200 130
rect 1080 51 1323 58
rect 1332 51 1440 58
<< metal6 >>
rect 1874 62 1882 593
rect 1890 2 1898 593
use logic  logic_0
timestamp 1575848640
transform 1 0 -327 0 1 504
box 87 2 327 70
use fadder  fadder_0
timestamp 1575778664
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1575848640
transform 1 0 -87 0 1 432
box 87 2 327 70
use fadder  fadder_1
timestamp 1575778664
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1575848640
transform 1 0 153 0 1 360
box 87 2 327 70
use fadder  fadder_2
timestamp 1575778664
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1575848640
transform 1 0 393 0 1 288
box 87 2 327 70
use fadder  fadder_3
timestamp 1575778664
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1575848640
transform 1 0 633 0 1 216
box 87 2 327 70
use fadder  fadder_4
timestamp 1575778664
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1575848640
transform 1 0 873 0 1 144
box 87 2 327 70
use fadder  fadder_5
timestamp 1575778664
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1575848640
transform 1 0 1113 0 1 72
box 87 2 327 70
use fadder  fadder_6
timestamp 1575778664
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1575778664
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1575848640
transform 1 0 1353 0 1 0
box 87 2 327 70
use mult  mult_0
timestamp 1575848640
transform 1 0 241 0 1 432
box -241 -432 1679 142
<< labels >>
rlabel metal6 1878 590 1878 590 5 Vdd
rlabel metal6 1894 589 1894 589 5 Gnd
<< end >>
