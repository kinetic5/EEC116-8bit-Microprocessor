magic
tech scmos
timestamp 1576011127
<< ntransistor >>
rect -47 4 -45 9
rect -27 4 -25 13
rect -17 4 -15 13
rect -7 4 -5 11
rect 3 4 5 11
rect 13 4 15 11
rect 23 4 25 11
rect 33 4 35 11
rect 43 4 45 11
rect 53 4 55 11
rect 63 4 65 11
rect 73 4 75 11
rect 83 4 85 11
rect 93 4 95 12
rect 103 4 105 12
rect 113 4 115 12
rect 123 4 125 12
rect 133 4 135 12
rect 143 4 145 12
rect 153 4 155 12
rect 163 4 165 12
rect 173 4 175 12
rect 183 4 185 12
rect 193 4 195 12
rect 203 4 205 12
rect 213 4 215 12
rect 223 4 225 12
rect 233 4 235 12
rect 243 4 245 12
rect 253 4 255 12
rect 263 4 265 12
rect 273 4 275 12
rect 283 4 285 12
rect 293 4 295 12
rect 303 4 305 12
rect 313 4 315 12
rect 323 4 325 12
rect 333 4 335 12
rect 343 4 345 12
rect 353 4 355 12
rect 363 4 365 12
rect 373 4 375 12
rect 383 4 385 12
<< ptransistor >>
rect -47 37 -45 47
rect -27 31 -25 47
rect -17 31 -15 47
rect -7 32 -5 47
rect 3 32 5 47
rect 13 32 15 47
rect 23 32 25 47
rect 33 32 35 47
rect 43 32 45 47
rect 53 32 55 47
rect 63 32 65 47
rect 73 32 75 47
rect 83 32 85 47
rect 93 31 95 47
rect 103 31 105 47
rect 113 31 115 47
rect 123 31 125 47
rect 133 31 135 47
rect 143 31 145 47
rect 153 31 155 47
rect 163 31 165 47
rect 173 31 175 47
rect 183 31 185 47
rect 193 31 195 47
rect 203 31 205 47
rect 213 31 215 47
rect 223 31 225 47
rect 233 31 235 47
rect 243 31 245 47
rect 253 31 255 47
rect 263 31 265 47
rect 273 31 275 47
rect 283 31 285 47
rect 293 31 295 47
rect 303 31 305 47
rect 313 31 315 47
rect 323 31 325 47
rect 333 31 335 47
rect 343 31 345 47
rect 353 31 355 47
rect 363 31 365 47
rect 373 31 375 47
rect 383 31 385 47
<< ndiffusion >>
rect -48 4 -47 9
rect -45 4 -44 9
rect -34 12 -27 13
rect -28 4 -27 12
rect -25 12 -17 13
rect -25 4 -24 12
rect -18 4 -17 12
rect -15 11 -8 13
rect 86 11 93 12
rect -15 4 -14 11
rect -8 4 -7 11
rect -5 4 -4 11
rect 2 4 3 11
rect 5 4 6 11
rect 12 4 13 11
rect 15 4 16 11
rect 22 4 23 11
rect 25 4 26 11
rect 32 4 33 11
rect 35 4 36 11
rect 42 4 43 11
rect 45 4 46 11
rect 52 4 53 11
rect 55 4 56 11
rect 62 4 63 11
rect 65 4 66 11
rect 72 4 73 11
rect 75 4 76 11
rect 82 4 83 11
rect 85 4 86 11
rect 92 4 93 11
rect 95 10 103 12
rect 95 4 96 10
rect 102 4 103 10
rect 105 11 113 12
rect 105 4 106 11
rect 112 4 113 11
rect 115 11 123 12
rect 115 4 116 11
rect 122 4 123 11
rect 125 11 133 12
rect 125 4 126 11
rect 132 4 133 11
rect 135 11 143 12
rect 135 4 136 11
rect 142 4 143 11
rect 145 11 153 12
rect 145 4 146 11
rect 152 4 153 11
rect 155 11 163 12
rect 155 4 156 11
rect 162 4 163 11
rect 165 11 173 12
rect 165 4 166 11
rect 172 4 173 11
rect 175 11 183 12
rect 175 4 176 11
rect 182 4 183 11
rect 185 11 193 12
rect 185 4 186 11
rect 192 4 193 11
rect 195 11 203 12
rect 195 4 196 11
rect 202 4 203 11
rect 205 11 213 12
rect 205 4 206 11
rect 212 4 213 11
rect 215 11 223 12
rect 215 4 216 11
rect 222 4 223 11
rect 225 11 233 12
rect 225 4 226 11
rect 232 4 233 11
rect 235 11 243 12
rect 235 4 236 11
rect 242 4 243 11
rect 245 11 253 12
rect 245 4 246 11
rect 252 4 253 11
rect 255 11 263 12
rect 255 4 256 11
rect 262 4 263 11
rect 265 11 273 12
rect 265 4 266 11
rect 272 4 273 11
rect 275 11 283 12
rect 275 4 276 11
rect 282 4 283 11
rect 285 11 293 12
rect 285 4 286 11
rect 292 4 293 11
rect 295 11 303 12
rect 295 4 296 11
rect 302 4 303 11
rect 305 11 313 12
rect 305 4 306 11
rect 312 4 313 11
rect 315 11 323 12
rect 315 4 316 11
rect 322 4 323 11
rect 325 11 333 12
rect 325 4 326 11
rect 332 4 333 11
rect 335 11 343 12
rect 335 4 336 11
rect 342 4 343 11
rect 345 11 353 12
rect 345 4 346 11
rect 352 4 353 11
rect 355 11 363 12
rect 355 4 356 11
rect 362 4 363 11
rect 365 11 373 12
rect 365 4 366 11
rect 372 4 373 11
rect 375 11 383 12
rect 375 4 376 11
rect 382 4 383 11
rect 385 11 392 12
rect 385 4 386 11
<< pdiffusion >>
rect -48 37 -47 47
rect -45 37 -44 47
rect -28 34 -27 47
rect -34 31 -27 34
rect -25 34 -24 47
rect -18 34 -17 47
rect -25 31 -17 34
rect -15 34 -14 47
rect -8 34 -7 47
rect -15 32 -7 34
rect -5 32 -4 47
rect 2 32 3 47
rect 5 32 6 47
rect 12 32 13 47
rect 15 32 16 47
rect 22 32 23 47
rect 25 32 26 47
rect 32 32 33 47
rect 35 32 36 47
rect 42 32 43 47
rect 45 32 46 47
rect 52 32 53 47
rect 55 32 56 47
rect 62 32 63 47
rect 65 32 66 47
rect 72 32 73 47
rect 75 32 76 47
rect 82 32 83 47
rect 85 32 86 47
rect 92 32 93 47
rect -15 31 -8 32
rect 86 31 93 32
rect 95 33 96 47
rect 102 33 103 47
rect 95 31 103 33
rect 105 32 106 47
rect 112 32 113 47
rect 105 31 113 32
rect 115 32 116 47
rect 122 32 123 47
rect 115 31 123 32
rect 125 32 126 47
rect 132 32 133 47
rect 125 31 133 32
rect 135 32 136 47
rect 142 32 143 47
rect 135 31 143 32
rect 145 32 146 47
rect 152 32 153 47
rect 145 31 153 32
rect 155 32 156 47
rect 162 32 163 47
rect 155 31 163 32
rect 165 32 166 47
rect 172 32 173 47
rect 165 31 173 32
rect 175 32 176 47
rect 182 32 183 47
rect 175 31 183 32
rect 185 32 186 47
rect 192 32 193 47
rect 185 31 193 32
rect 195 32 196 47
rect 202 32 203 47
rect 195 31 203 32
rect 205 32 206 47
rect 212 32 213 47
rect 205 31 213 32
rect 215 32 216 47
rect 222 32 223 47
rect 215 31 223 32
rect 225 32 226 47
rect 232 32 233 47
rect 225 31 233 32
rect 235 32 236 47
rect 242 32 243 47
rect 235 31 243 32
rect 245 32 246 47
rect 252 32 253 47
rect 245 31 253 32
rect 255 32 256 47
rect 262 32 263 47
rect 255 31 263 32
rect 265 32 266 47
rect 272 32 273 47
rect 265 31 273 32
rect 275 32 276 47
rect 282 32 283 47
rect 275 31 283 32
rect 285 32 286 47
rect 292 32 293 47
rect 285 31 293 32
rect 295 32 296 47
rect 302 32 303 47
rect 295 31 303 32
rect 305 32 306 47
rect 312 32 313 47
rect 305 31 313 32
rect 315 32 316 47
rect 322 32 323 47
rect 315 31 323 32
rect 325 32 326 47
rect 332 32 333 47
rect 325 31 333 32
rect 335 32 336 47
rect 342 32 343 47
rect 335 31 343 32
rect 345 32 346 47
rect 352 32 353 47
rect 345 31 353 32
rect 355 32 356 47
rect 362 32 363 47
rect 355 31 363 32
rect 365 32 366 47
rect 372 32 373 47
rect 365 31 373 32
rect 375 32 376 47
rect 382 32 383 47
rect 375 31 383 32
rect 385 32 386 47
rect 385 31 390 32
<< ndcontact >>
rect -54 4 -48 9
rect -44 4 -38 9
rect -34 4 -28 12
rect -14 4 -8 11
rect 6 4 12 11
rect 26 4 32 11
rect 46 4 52 11
rect 66 4 72 11
rect 86 4 92 11
rect 106 3 112 11
rect 126 3 132 11
rect 146 3 152 11
rect 166 3 172 11
rect 186 3 192 11
rect 206 3 212 11
rect 226 3 232 11
rect 246 3 252 11
rect 266 3 272 11
rect 286 3 292 11
rect 306 3 312 11
rect 326 3 332 11
rect 346 3 352 11
rect 366 3 372 11
rect 386 3 392 11
<< pdcontact >>
rect -54 37 -48 47
rect -44 37 -38 47
rect -34 34 -28 47
rect -14 34 -8 47
rect 6 32 12 47
rect 26 32 32 47
rect 46 32 52 47
rect 66 32 72 47
rect 86 32 92 47
rect 106 32 112 47
rect 126 32 132 47
rect 146 32 152 47
rect 166 32 172 47
rect 186 32 192 47
rect 206 32 212 47
rect 226 32 232 47
rect 246 32 252 47
rect 266 32 272 47
rect 286 32 292 47
rect 306 32 312 47
rect 326 32 332 47
rect 346 32 352 47
rect 366 32 372 47
rect 386 32 392 47
<< polysilicon >>
rect -57 1 -55 50
rect -47 47 -45 50
rect -47 33 -45 37
rect -47 9 -45 12
rect -47 1 -45 4
rect -37 1 -35 50
rect -27 47 -25 50
rect -17 47 -15 50
rect -7 47 -5 50
rect 3 47 5 50
rect 13 47 15 50
rect 23 47 25 50
rect 33 47 35 50
rect 43 47 45 50
rect 53 47 55 50
rect 63 47 65 50
rect 73 47 75 50
rect 83 47 85 50
rect 93 47 95 50
rect -27 28 -25 31
rect -17 28 -15 31
rect -7 28 -5 32
rect 3 29 5 32
rect 13 29 15 32
rect 23 29 25 32
rect 33 29 35 32
rect 43 29 45 32
rect 53 29 55 32
rect 63 29 65 32
rect 73 29 75 32
rect 83 29 85 32
rect 103 47 105 50
rect 113 47 115 50
rect 123 47 125 50
rect 133 47 135 50
rect 143 47 145 50
rect 153 47 155 50
rect 163 47 165 50
rect 173 47 175 50
rect 183 47 185 50
rect 193 47 195 50
rect 203 47 205 50
rect 213 47 215 50
rect 223 47 225 50
rect 233 47 235 50
rect 243 47 245 50
rect 253 47 255 50
rect 263 47 265 50
rect 273 47 275 50
rect 283 47 285 50
rect 293 47 295 50
rect 303 47 305 50
rect 313 47 315 50
rect 323 47 325 50
rect 333 47 335 50
rect 343 47 345 50
rect 353 47 355 50
rect 363 47 365 50
rect 373 47 375 50
rect 383 47 385 50
rect 93 29 95 31
rect 103 29 105 31
rect 113 29 115 31
rect 123 29 125 31
rect 133 29 135 31
rect 143 29 145 31
rect 153 29 155 31
rect 163 29 165 31
rect 173 29 175 31
rect 183 29 185 31
rect 193 29 195 31
rect 203 29 205 31
rect 213 29 215 31
rect 223 29 225 31
rect 233 29 235 31
rect 243 29 245 31
rect 253 29 255 31
rect 263 29 265 31
rect 273 29 275 31
rect 283 29 285 31
rect 293 29 295 31
rect 303 29 305 31
rect 313 29 315 31
rect 323 29 325 31
rect 333 29 335 31
rect 343 29 345 31
rect 353 29 355 31
rect 363 29 365 31
rect 373 29 375 31
rect 383 29 385 31
rect -27 13 -25 15
rect -17 13 -15 15
rect -7 11 -5 15
rect 3 11 5 14
rect 13 11 15 14
rect 23 11 25 14
rect 33 11 35 14
rect 43 11 45 14
rect 53 11 55 14
rect 63 11 65 14
rect 73 11 75 14
rect 83 11 85 14
rect 93 12 95 14
rect 103 12 105 14
rect 113 12 115 14
rect 123 12 125 14
rect 133 12 135 14
rect 143 12 145 14
rect 153 12 155 14
rect 163 12 165 14
rect 173 12 175 14
rect 183 12 185 14
rect 193 12 195 14
rect 203 12 205 14
rect 213 12 215 14
rect 223 12 225 14
rect 233 12 235 14
rect 243 12 245 14
rect 253 12 255 14
rect 263 12 265 14
rect 273 12 275 14
rect 283 12 285 14
rect 293 12 295 14
rect 303 12 305 14
rect 313 12 315 14
rect 323 12 325 14
rect 333 12 335 14
rect 343 12 345 14
rect 353 12 355 14
rect 363 12 365 14
rect 373 12 375 14
rect 383 12 385 14
rect -27 1 -25 4
rect -17 1 -15 4
rect -7 1 -5 4
rect 3 1 5 4
rect 13 1 15 4
rect 23 1 25 4
rect 33 1 35 4
rect 43 1 45 4
rect 53 1 55 4
rect 63 1 65 4
rect 73 1 75 4
rect 83 1 85 4
rect 93 1 95 4
rect 103 1 105 4
rect 113 1 115 4
rect 123 1 125 4
rect 133 1 135 4
rect 143 1 145 4
rect 153 1 155 4
rect 163 1 165 4
rect 173 1 175 4
rect 183 1 185 4
rect 193 1 195 4
rect 203 1 205 4
rect 213 1 215 4
rect 223 1 225 4
rect 233 1 235 4
rect 243 1 245 4
rect 253 1 255 4
rect 263 1 265 4
rect 273 1 275 4
rect 283 1 285 4
rect 293 1 295 4
rect 303 1 305 4
rect 313 1 315 4
rect 323 1 325 4
rect 333 1 335 4
rect 343 1 345 4
rect 353 1 355 4
rect 363 1 365 4
rect 373 1 375 4
rect 383 1 385 4
rect 393 1 395 50
rect 403 1 405 50
<< polycontact >>
rect -29 15 -23 28
rect -19 15 -13 28
rect 1 14 7 29
rect 11 14 17 29
rect 21 14 27 29
rect 31 14 37 29
rect 41 14 47 29
rect 51 14 57 29
rect 61 14 67 29
rect 71 14 77 29
rect 81 14 87 29
rect 101 14 107 29
rect 111 14 117 29
rect 121 14 127 29
rect 131 14 137 29
rect 141 14 147 29
rect 151 14 157 29
rect 161 14 167 29
rect 171 14 177 29
rect 181 14 187 29
rect 191 14 197 29
rect 201 14 207 29
rect 211 14 217 29
rect 221 14 227 29
rect 231 14 237 29
rect 241 14 247 29
rect 251 14 257 29
rect 261 14 267 29
rect 271 14 277 29
rect 281 14 287 29
rect 291 14 297 29
rect 301 14 307 29
rect 311 14 317 29
rect 321 14 327 29
rect 331 14 337 29
rect 341 14 347 29
rect 351 14 357 29
rect 361 14 367 29
rect 371 14 377 29
rect 381 14 387 29
<< metal1 >>
rect -61 51 409 59
rect -54 47 -48 51
rect -34 47 -28 51
rect -14 47 -8 51
rect 6 47 12 51
rect 26 47 32 51
rect 46 47 52 51
rect 66 47 72 51
rect 86 47 92 51
rect -38 37 -37 47
rect -41 31 -37 37
rect 106 47 112 51
rect 126 47 132 51
rect 146 47 152 51
rect 166 47 172 51
rect 186 47 192 51
rect 206 47 212 51
rect 226 47 232 51
rect 246 47 252 51
rect 266 47 272 51
rect 286 47 292 51
rect 306 47 312 51
rect 326 47 332 51
rect 346 47 352 51
rect 366 47 372 51
rect 386 47 392 51
rect -41 28 -16 31
rect -9 28 1 29
rect -41 15 -29 28
rect -23 15 -19 28
rect -3 15 1 28
rect -41 9 -37 15
rect -9 14 1 15
rect 7 14 11 29
rect 17 14 21 29
rect 27 14 31 29
rect 37 14 41 29
rect 47 14 51 29
rect 57 14 61 29
rect 67 14 71 29
rect 77 14 81 29
rect 97 14 101 29
rect 107 14 111 29
rect 117 14 121 29
rect 127 14 131 29
rect 137 14 141 29
rect 147 14 151 29
rect 157 14 161 29
rect 167 14 171 29
rect 177 14 181 29
rect 187 14 191 29
rect 197 14 201 29
rect 207 14 211 29
rect 217 14 221 29
rect 227 14 231 29
rect 237 14 241 29
rect 247 14 251 29
rect 257 14 261 29
rect 267 14 271 29
rect 277 14 281 29
rect 287 14 291 29
rect 297 14 301 29
rect 307 14 311 29
rect 317 14 321 29
rect 327 14 331 29
rect 337 14 341 29
rect 347 14 351 29
rect 357 14 361 29
rect 367 14 371 29
rect 377 14 381 29
rect -38 4 -37 9
rect -54 -1 -48 4
rect -34 -1 -28 4
rect -14 -1 -8 4
rect 6 -1 12 4
rect 26 -1 32 4
rect 46 -1 52 4
rect 66 -1 72 4
rect 86 -1 92 4
rect 106 -1 112 3
rect 126 -1 132 3
rect 146 -1 152 3
rect 166 -1 172 3
rect 186 -1 192 3
rect 206 -1 212 3
rect 226 -1 232 3
rect 246 -1 252 3
rect 266 -1 272 3
rect 286 -1 292 3
rect 306 -1 312 3
rect 326 -1 332 3
rect 346 -1 352 3
rect 366 -1 372 3
rect 386 -1 392 3
rect -61 -9 409 -1
<< pm12contact >>
rect -49 12 -44 33
rect -9 15 -3 28
rect 91 14 97 29
<< pdm12contact >>
rect -24 34 -18 47
rect -4 32 2 47
rect 16 32 22 47
rect 36 32 42 47
rect 56 32 62 47
rect 76 32 82 47
rect 96 33 102 48
rect 116 32 122 48
rect 136 32 142 48
rect 156 32 162 48
rect 176 32 182 48
rect 196 32 202 48
rect 216 32 222 48
rect 236 32 242 48
rect 256 32 262 48
rect 276 32 282 48
rect 296 32 302 48
rect 316 32 322 48
rect 336 32 342 48
rect 356 32 362 48
rect 376 32 382 48
<< ndm12contact >>
rect -24 4 -18 12
rect -4 2 2 11
rect 16 2 22 11
rect 36 2 42 11
rect 56 2 62 11
rect 76 2 82 11
rect 96 2 102 10
rect 116 2 122 11
rect 136 2 142 11
rect 156 2 162 11
rect 176 2 182 11
rect 196 2 202 11
rect 216 2 222 11
rect 236 2 242 11
rect 256 2 262 11
rect 276 2 282 11
rect 296 2 302 11
rect 316 2 322 11
rect 336 2 342 11
rect 356 2 362 11
rect 376 2 382 11
<< metal2 >>
rect -18 34 -14 47
rect -24 28 -14 34
rect 2 32 16 47
rect 22 32 36 47
rect 42 32 56 47
rect 62 32 76 47
rect 102 33 116 48
rect 16 29 82 32
rect 101 32 116 33
rect 122 32 136 48
rect 142 32 156 48
rect 162 32 176 48
rect 182 32 196 48
rect 202 32 216 48
rect 222 32 236 48
rect 242 32 256 48
rect 262 32 276 48
rect 282 32 296 48
rect 302 32 316 48
rect 322 32 336 48
rect 342 32 356 48
rect 362 32 376 48
rect 382 36 390 48
rect 382 32 388 36
rect -24 15 -9 28
rect -24 12 -14 15
rect -18 4 -14 12
rect 16 14 91 29
rect 16 11 82 14
rect 2 2 16 11
rect 22 2 36 11
rect 42 2 56 11
rect 62 2 76 11
rect 101 12 388 32
rect 101 11 390 12
rect 101 10 116 11
rect 102 2 116 10
rect 122 2 136 11
rect 142 2 156 11
rect 162 2 176 11
rect 182 2 196 11
rect 202 2 216 11
rect 222 2 236 11
rect 242 2 256 11
rect 262 2 276 11
rect 282 2 296 11
rect 302 2 316 11
rect 322 2 336 11
rect 342 2 356 11
rect 362 2 376 11
rect 382 2 390 11
<< m3contact >>
rect -54 12 -49 33
rect 388 12 402 36
<< labels >>
rlabel m3contact -53 21 -53 21 3 in
rlabel m3contact 399 23 399 23 1 out
rlabel metal1 -51 -6 -51 -6 1 Gnd
rlabel metal1 -50 54 -50 54 5 Vdd
<< end >>
