magic
tech scmos
timestamp 1575778145
<< error_s >>
rect 308 445 318 446
rect 548 373 558 374
rect 788 301 798 302
rect 1028 229 1038 230
rect 1268 157 1278 158
rect 1508 85 1518 86
rect 1748 13 1758 14
<< metal6 >>
rect 1874 62 1882 593
rect 1890 2 1898 593
use logic  logic_0
timestamp 1575777673
transform 1 0 -327 0 1 504
box 87 2 327 70
use fadder  fadder_0
timestamp 1575777673
transform 1 0 -156 0 1 430
box -24 4 156 72
use logic  logic_1
timestamp 1575777673
transform 1 0 -87 0 1 432
box 87 2 327 70
use fadder  fadder_1
timestamp 1575777673
transform 1 0 84 0 1 358
box -24 4 156 72
use logic  logic_2
timestamp 1575777673
transform 1 0 153 0 1 360
box 87 2 327 70
use fadder  fadder_2
timestamp 1575777673
transform 1 0 324 0 1 286
box -24 4 156 72
use logic  logic_3
timestamp 1575777673
transform 1 0 393 0 1 288
box 87 2 327 70
use fadder  fadder_3
timestamp 1575777673
transform 1 0 564 0 1 214
box -24 4 156 72
use logic  logic_4
timestamp 1575777673
transform 1 0 633 0 1 216
box 87 2 327 70
use fadder  fadder_4
timestamp 1575777673
transform 1 0 804 0 1 142
box -24 4 156 72
use logic  logic_5
timestamp 1575777673
transform 1 0 873 0 1 144
box 87 2 327 70
use fadder  fadder_5
timestamp 1575777673
transform 1 0 1044 0 1 70
box -24 4 156 72
use logic  logic_6
timestamp 1575777673
transform 1 0 1113 0 1 72
box 87 2 327 70
use fadder  fadder_6
timestamp 1575777673
transform 1 0 1104 0 1 -2
box -24 4 156 72
use fadder  fadder_7
timestamp 1575777673
transform 1 0 1284 0 1 -2
box -24 4 156 72
use logic  logic_7
timestamp 1575777673
transform 1 0 1353 0 1 0
box 87 2 327 70
use mult  mult_0
timestamp 1575778145
transform 1 0 241 0 1 432
box -241 -432 1679 142
<< labels >>
rlabel metal6 1878 590 1878 590 5 Vdd
rlabel metal6 1894 589 1894 589 5 Gnd
<< end >>
