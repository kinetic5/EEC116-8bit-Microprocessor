magic
tech scmos
timestamp 1575938163
<< ntransistor >>
rect -62 -97 -60 -93
rect -52 -97 -50 -93
rect -42 -97 -40 -93
rect -32 -97 -30 -93
rect -12 -97 -10 -93
rect -2 -97 0 -93
rect 8 -97 10 -93
rect 18 -97 20 -93
rect -22 -105 -20 -101
rect 38 -97 40 -93
rect 28 -105 30 -101
rect 76 -99 78 -93
rect 86 -97 88 -93
rect 66 -108 68 -104
rect 106 -101 108 -93
rect 116 -101 118 -93
<< ptransistor >>
rect -22 -71 -20 -65
rect -62 -81 -60 -75
rect -52 -81 -50 -75
rect -42 -81 -40 -75
rect -32 -81 -30 -75
rect 28 -71 30 -65
rect -12 -81 -10 -75
rect -2 -81 0 -75
rect 8 -81 10 -75
rect 18 -81 20 -75
rect 38 -81 40 -75
rect 66 -70 68 -64
rect 76 -81 78 -75
rect 86 -81 88 -75
rect 106 -81 108 -69
rect 116 -81 118 -69
<< ndiffusion >>
rect -63 -97 -62 -93
rect -60 -97 -59 -93
rect -53 -97 -52 -93
rect -50 -97 -49 -93
rect -43 -97 -42 -93
rect -40 -97 -39 -93
rect -33 -97 -32 -93
rect -30 -97 -29 -93
rect -13 -97 -12 -93
rect -10 -97 -9 -93
rect -3 -97 -2 -93
rect 0 -97 1 -93
rect 7 -97 8 -93
rect 10 -97 11 -93
rect 17 -97 18 -93
rect 20 -97 21 -93
rect -19 -101 -14 -97
rect -27 -105 -22 -101
rect -20 -105 -14 -101
rect -27 -109 -23 -105
rect 37 -97 38 -93
rect 40 -97 47 -93
rect 23 -105 28 -101
rect 30 -105 31 -101
rect 23 -109 27 -105
rect 41 -102 47 -97
rect 69 -95 76 -93
rect 69 -99 70 -95
rect 75 -99 76 -95
rect 78 -97 80 -93
rect 85 -97 86 -93
rect 88 -97 89 -93
rect 78 -99 82 -97
rect 64 -105 66 -104
rect 59 -108 66 -105
rect 68 -108 74 -104
rect 69 -112 74 -108
rect 105 -101 106 -93
rect 108 -101 109 -93
rect 115 -101 116 -93
rect 118 -101 119 -93
<< pdiffusion >>
rect -23 -71 -22 -65
rect -20 -71 -14 -65
rect -63 -81 -62 -75
rect -60 -81 -59 -75
rect -53 -81 -52 -75
rect -50 -81 -49 -75
rect -43 -81 -42 -75
rect -40 -81 -39 -75
rect -33 -81 -32 -75
rect -30 -81 -29 -75
rect -19 -75 -14 -71
rect 27 -71 28 -65
rect 30 -70 31 -65
rect 30 -71 37 -70
rect -13 -81 -12 -75
rect -10 -81 -9 -75
rect -3 -81 -2 -75
rect 0 -81 1 -75
rect 7 -81 8 -75
rect 10 -81 11 -75
rect 17 -81 18 -75
rect 20 -81 21 -75
rect 41 -75 47 -72
rect 37 -81 38 -75
rect 40 -81 47 -75
rect 69 -64 74 -60
rect 65 -70 66 -64
rect 68 -70 74 -64
rect 69 -80 71 -75
rect 75 -80 76 -75
rect 69 -81 76 -80
rect 78 -81 80 -75
rect 85 -81 86 -75
rect 88 -81 89 -75
rect 105 -81 106 -69
rect 108 -81 109 -69
rect 115 -81 116 -69
rect 118 -81 119 -69
<< ndcontact >>
rect -69 -97 -63 -93
rect -59 -97 -53 -93
rect -49 -97 -43 -93
rect -39 -97 -33 -93
rect -29 -97 -23 -93
rect -19 -97 -13 -93
rect -9 -97 -3 -93
rect 1 -97 7 -93
rect 11 -97 17 -93
rect 21 -97 26 -93
rect 31 -97 37 -93
rect 41 -107 47 -102
rect -27 -113 -23 -109
rect 23 -113 27 -109
rect 59 -105 64 -101
rect 70 -99 75 -95
rect 80 -97 85 -93
rect 99 -101 105 -93
rect 119 -101 125 -93
rect 69 -116 74 -112
<< pdcontact >>
rect 69 -60 75 -56
rect -29 -71 -23 -65
rect -69 -81 -63 -75
rect -59 -81 -53 -75
rect -49 -81 -43 -75
rect -39 -81 -33 -75
rect -29 -81 -23 -75
rect 21 -71 27 -65
rect -19 -81 -13 -75
rect -9 -81 -3 -75
rect 1 -81 7 -75
rect 11 -81 17 -75
rect 21 -81 26 -75
rect 41 -72 47 -67
rect 31 -81 37 -75
rect 59 -70 65 -64
rect 71 -80 75 -75
rect 80 -81 85 -75
rect 99 -81 105 -69
rect 119 -81 125 -69
<< polysilicon >>
rect -72 -109 -70 -63
rect -62 -65 -60 -63
rect -52 -65 -50 -63
rect -62 -75 -60 -71
rect -52 -75 -50 -71
rect -42 -75 -40 -63
rect -32 -75 -30 -63
rect -22 -65 -20 -62
rect -12 -65 -10 -63
rect -2 -65 0 -63
rect -62 -84 -60 -81
rect -52 -84 -50 -81
rect -42 -84 -40 -81
rect -62 -93 -60 -90
rect -52 -93 -50 -90
rect -42 -93 -40 -90
rect -32 -93 -30 -81
rect -22 -84 -20 -71
rect -12 -75 -10 -71
rect -2 -75 0 -71
rect 8 -75 10 -63
rect 18 -75 20 -63
rect 28 -65 30 -62
rect -12 -84 -10 -81
rect -2 -84 0 -81
rect 8 -84 10 -81
rect -62 -101 -60 -97
rect -52 -101 -50 -97
rect -62 -109 -60 -107
rect -52 -109 -50 -107
rect -42 -109 -40 -97
rect -32 -100 -30 -97
rect -22 -101 -20 -90
rect -12 -93 -10 -90
rect -2 -93 0 -90
rect 8 -93 10 -90
rect 18 -93 20 -81
rect 28 -84 30 -71
rect 38 -75 40 -63
rect 38 -84 40 -81
rect -12 -101 -10 -97
rect -2 -101 0 -97
rect -32 -109 -30 -105
rect -22 -109 -20 -105
rect -12 -109 -10 -107
rect -2 -108 0 -107
rect 8 -108 10 -97
rect 18 -100 20 -97
rect 28 -101 30 -90
rect 38 -93 40 -90
rect 18 -108 20 -105
rect 28 -108 30 -105
rect 38 -108 40 -97
rect 48 -110 50 -63
rect 56 -110 58 -62
rect 66 -64 68 -61
rect 76 -67 78 -62
rect 86 -66 88 -62
rect 66 -80 68 -70
rect 76 -75 78 -72
rect 86 -75 88 -71
rect 76 -84 78 -81
rect 86 -84 88 -81
rect 66 -88 68 -84
rect 66 -104 68 -92
rect 76 -93 78 -90
rect 86 -93 88 -90
rect 76 -102 78 -99
rect 86 -103 88 -97
rect 66 -111 68 -108
rect 76 -110 78 -107
rect 86 -110 88 -108
rect 96 -110 98 -62
rect 106 -69 108 -62
rect 116 -69 118 -62
rect 106 -84 108 -81
rect 116 -84 118 -81
rect 106 -93 108 -90
rect 116 -93 118 -90
rect 106 -110 108 -101
rect 116 -110 118 -101
rect 126 -110 128 -62
<< polycontact >>
rect -42 -90 -38 -84
rect -24 -90 -20 -84
rect 8 -90 12 -84
rect 28 -90 32 -84
rect 64 -84 68 -80
rect 104 -90 110 -84
rect 114 -90 120 -84
<< metal1 >>
rect -76 -56 132 -52
rect -76 -60 69 -56
rect 75 -60 132 -56
rect -39 -75 -33 -60
rect -29 -65 -23 -60
rect 11 -75 17 -60
rect 21 -65 27 -60
rect 41 -67 47 -60
rect 54 -70 59 -64
rect 65 -70 66 -64
rect -69 -83 -63 -81
rect -69 -93 -63 -91
rect -59 -88 -53 -81
rect -50 -81 -49 -75
rect -50 -93 -45 -81
rect -29 -84 -23 -81
rect -38 -90 -24 -84
rect -29 -93 -23 -90
rect -17 -93 -13 -81
rect -50 -97 -49 -93
rect -40 -97 -39 -93
rect -9 -86 -3 -81
rect -9 -93 -3 -91
rect 0 -81 1 -75
rect 29 -81 31 -75
rect 37 -80 41 -75
rect 37 -81 47 -80
rect 0 -93 5 -81
rect 21 -84 25 -81
rect 29 -84 33 -81
rect 12 -90 18 -84
rect 32 -90 33 -84
rect 21 -93 25 -90
rect 29 -93 33 -90
rect 0 -97 1 -93
rect 10 -97 11 -93
rect 29 -97 31 -93
rect 37 -94 47 -93
rect 37 -97 41 -94
rect -40 -112 -36 -97
rect -76 -113 -27 -112
rect 10 -112 14 -97
rect 29 -98 41 -97
rect 54 -94 60 -70
rect 99 -69 105 -60
rect 119 -69 125 -60
rect 75 -80 77 -75
rect 59 -99 60 -94
rect 75 -99 77 -95
rect 80 -84 85 -81
rect 80 -90 104 -84
rect 110 -90 114 -84
rect 80 -93 85 -90
rect 54 -101 60 -99
rect 54 -105 59 -101
rect -23 -113 23 -112
rect 41 -112 47 -107
rect 99 -112 105 -101
rect 119 -112 125 -101
rect 27 -113 69 -112
rect -76 -116 69 -113
rect 74 -116 132 -112
rect -76 -120 132 -116
<< pm12contact >>
rect -63 -71 -58 -65
rect -54 -71 -49 -65
rect -13 -71 -8 -65
rect -4 -71 1 -65
rect 36 -90 42 -84
rect -63 -107 -58 -101
rect -54 -107 -49 -101
rect -33 -105 -28 -100
rect -13 -107 -8 -101
rect -4 -107 1 -101
rect 75 -72 80 -67
rect 84 -71 89 -66
rect 17 -105 22 -100
rect 75 -107 80 -102
rect 84 -108 89 -103
<< pdm12contact >>
rect 31 -70 37 -65
rect 89 -81 95 -75
rect 109 -81 115 -69
<< ndm12contact >>
rect 89 -99 95 -93
rect 109 -101 115 -93
rect 31 -106 37 -101
<< metal2 >>
rect -64 -61 37 -55
rect -64 -65 -58 -61
rect -4 -65 2 -61
rect -64 -71 -63 -65
rect 1 -71 2 -65
rect 7 -65 37 -61
rect -33 -100 -28 -98
rect -49 -107 -48 -101
rect -54 -111 -48 -107
rect -14 -107 -13 -101
rect -14 -111 -8 -107
rect 7 -111 13 -65
rect 54 -71 75 -66
rect 27 -80 36 -74
rect 30 -90 36 -80
rect 54 -94 59 -71
rect 72 -72 75 -71
rect 17 -100 22 -99
rect 31 -111 37 -106
rect 63 -102 68 -80
rect 89 -87 95 -81
rect 89 -93 105 -87
rect 63 -107 75 -102
rect -63 -117 37 -111
rect 99 -112 105 -93
<< m3contact >>
rect -49 -71 -43 -65
rect -19 -71 -13 -65
rect -33 -98 -28 -93
rect -69 -107 -63 -101
rect -4 -101 2 -96
rect 19 -80 27 -72
rect 89 -71 94 -66
rect 17 -99 22 -94
rect 89 -108 94 -103
rect 109 -93 119 -81
<< m123contact >>
rect -69 -91 -63 -83
rect -59 -93 -53 -88
rect -9 -91 -3 -86
rect 41 -80 47 -75
rect 18 -90 25 -84
rect 41 -99 47 -94
rect 54 -99 59 -94
rect 63 -80 68 -75
rect 72 -95 77 -80
<< metal3 >>
rect -49 -61 47 -55
rect -49 -65 -43 -61
rect -19 -65 -13 -61
rect 41 -75 47 -61
rect 63 -71 89 -66
rect 63 -75 68 -71
rect -9 -86 14 -83
rect -3 -88 14 -86
rect -59 -97 -33 -93
rect 9 -94 14 -88
rect 25 -90 72 -84
rect 9 -98 17 -94
rect 11 -99 17 -98
rect -4 -103 2 -101
rect 41 -103 47 -99
rect -63 -107 47 -103
rect -69 -109 47 -107
rect 54 -103 59 -99
rect 54 -108 89 -103
<< labels >>
rlabel m123contact -66 -87 -66 -87 1 d
rlabel m123contact -6 -88 -6 -88 1 transm23_out
rlabel metal1 -56 -86 -56 -86 1 transm01_out
rlabel pdm12contact 34 -68 34 -68 1 _clk
rlabel m3contact 23 -73 23 -73 1 clk
rlabel metal1 -71 -56 -71 -56 4 Vdd
rlabel metal1 -72 -115 -72 -115 2 Gnd
rlabel metal1 31 -92 31 -92 1 _nclk
rlabel metal3 48 -87 48 -87 1 nq
rlabel metal2 92 -86 92 -86 1 D
rlabel metal1 82 -88 82 -88 1 mux_out
rlabel metal1 80 -116 80 -116 1 Gnd
rlabel metal1 116 -56 116 -56 7 Vdd
rlabel m123contact 65 -78 65 -78 1 enable
rlabel m3contact 113 -88 113 -88 1 Q
<< end >>
