magic
tech scmos
timestamp 1575836395
<< error_s >>
rect 294 21 295 22
<< ntransistor >>
rect 301 21 303 33
rect 311 21 313 33
rect 331 32 333 36
rect 321 21 323 27
rect 341 29 343 33
rect 371 29 373 33
rect 381 29 383 33
rect 391 29 393 33
rect 401 29 403 33
rect 361 21 363 25
rect 431 29 433 33
rect 441 29 443 33
rect 461 29 463 33
rect 471 29 473 33
rect 421 21 423 25
<< ptransistor >>
rect 301 49 303 67
rect 311 49 313 67
rect 321 59 323 67
rect 331 49 333 55
rect 341 53 343 59
rect 361 62 363 67
rect 371 53 373 59
rect 381 53 383 59
rect 391 53 393 59
rect 401 53 403 59
rect 421 62 423 67
rect 431 53 433 59
rect 441 53 443 59
rect 461 53 463 59
rect 471 53 473 59
<< ndiffusion >>
rect 300 21 301 33
rect 303 32 311 33
rect 303 21 304 32
rect 310 21 311 32
rect 313 21 314 33
rect 329 32 331 36
rect 333 32 334 36
rect 320 21 321 27
rect 323 21 324 27
rect 340 29 341 33
rect 343 29 345 33
rect 369 29 371 33
rect 373 29 374 33
rect 380 29 381 33
rect 383 29 385 33
rect 389 29 391 33
rect 393 29 394 33
rect 399 29 401 33
rect 403 29 404 33
rect 408 29 409 33
rect 359 21 361 25
rect 363 21 368 25
rect 430 29 431 33
rect 433 29 435 33
rect 439 29 441 33
rect 443 29 444 33
rect 460 29 461 33
rect 463 29 464 33
rect 470 29 471 33
rect 473 29 474 33
rect 418 21 421 25
rect 423 21 429 25
rect 364 18 368 21
rect 424 18 428 21
<< pdiffusion >>
rect 300 50 301 67
rect 294 49 301 50
rect 303 50 304 67
rect 310 50 311 67
rect 303 49 311 50
rect 313 50 314 67
rect 320 59 321 67
rect 323 59 324 67
rect 313 49 320 50
rect 330 49 331 55
rect 333 53 334 55
rect 340 53 341 59
rect 343 53 345 59
rect 333 49 340 53
rect 364 67 368 70
rect 424 67 428 71
rect 359 62 361 67
rect 363 62 368 67
rect 365 58 371 59
rect 369 53 371 58
rect 373 53 374 59
rect 380 53 381 59
rect 383 53 384 59
rect 390 53 391 59
rect 393 53 394 59
rect 400 53 401 59
rect 403 53 404 59
rect 408 53 409 59
rect 419 62 421 67
rect 423 62 428 67
rect 425 58 431 59
rect 429 53 431 58
rect 433 53 435 59
rect 439 53 441 59
rect 443 58 449 59
rect 443 53 444 58
rect 460 53 461 59
rect 463 53 464 59
rect 470 53 471 59
rect 473 54 474 59
rect 473 53 479 54
<< ndcontact >>
rect 294 21 300 33
rect 314 21 320 33
rect 325 32 329 36
rect 334 29 340 36
rect 345 29 349 33
rect 365 29 369 33
rect 374 29 380 33
rect 385 29 389 33
rect 394 29 399 33
rect 404 29 408 33
rect 355 21 359 25
rect 426 29 430 33
rect 435 29 439 33
rect 444 29 450 33
rect 455 29 460 33
rect 464 29 470 33
rect 474 29 479 33
rect 414 21 418 25
rect 364 14 368 18
rect 424 14 428 18
<< pdcontact >>
rect 364 70 368 74
rect 424 71 428 75
rect 294 50 300 67
rect 314 50 320 67
rect 324 49 330 55
rect 334 53 340 59
rect 345 53 349 59
rect 355 62 359 67
rect 365 53 369 58
rect 374 53 380 59
rect 384 53 390 59
rect 394 53 400 59
rect 404 53 408 59
rect 415 62 419 67
rect 425 53 429 58
rect 435 53 439 59
rect 455 53 460 59
rect 464 53 470 59
rect 474 54 479 59
<< psubstratepcontact >>
rect 334 11 350 18
rect 388 11 400 18
rect 434 12 442 18
<< nsubstratencontact >>
rect 388 70 403 77
rect 432 71 441 77
<< polysilicon >>
rect 301 67 303 70
rect 311 67 313 70
rect 321 67 323 70
rect 301 46 303 49
rect 311 46 313 49
rect 321 47 323 59
rect 331 55 333 70
rect 341 59 343 70
rect 331 44 333 49
rect 341 44 343 53
rect 301 33 303 36
rect 311 33 313 36
rect 321 27 323 38
rect 331 36 333 39
rect 331 21 333 32
rect 341 33 343 39
rect 341 21 343 29
rect 351 21 353 70
rect 361 67 363 70
rect 421 67 423 70
rect 361 41 363 62
rect 371 59 373 62
rect 381 59 383 62
rect 391 59 393 67
rect 401 59 403 67
rect 371 46 373 53
rect 381 46 383 53
rect 391 41 393 53
rect 361 25 363 36
rect 371 33 373 40
rect 381 33 383 40
rect 391 33 393 36
rect 401 33 403 53
rect 371 26 373 29
rect 381 26 383 29
rect 391 21 393 29
rect 401 26 403 29
rect 411 21 413 67
rect 421 41 423 62
rect 431 59 433 62
rect 441 59 443 62
rect 431 46 433 53
rect 441 46 443 53
rect 421 25 423 36
rect 431 33 433 40
rect 441 33 443 40
rect 431 26 433 29
rect 441 26 443 29
rect 451 26 453 62
rect 461 59 463 62
rect 471 59 473 62
rect 461 50 463 53
rect 461 33 463 45
rect 471 41 473 53
rect 471 33 473 36
rect 461 26 463 29
rect 471 26 473 29
rect 481 26 483 62
rect 301 18 303 21
rect 311 18 313 21
rect 321 18 323 21
rect 361 18 363 21
rect 421 18 423 21
<< polycontact >>
rect 321 38 325 47
rect 330 39 334 44
rect 469 36 473 41
<< metal1 >>
rect 247 77 487 78
rect 247 74 388 77
rect 247 70 364 74
rect 368 70 388 74
rect 403 75 432 77
rect 403 71 424 75
rect 428 71 432 75
rect 441 71 487 77
rect 403 70 487 71
rect 294 67 300 70
rect 314 67 320 70
rect 334 59 340 70
rect 354 62 355 67
rect 323 49 324 55
rect 323 47 327 49
rect 325 38 327 47
rect 334 39 338 44
rect 323 36 327 38
rect 323 32 325 36
rect 346 33 350 48
rect 349 29 350 33
rect 354 32 357 62
rect 394 59 400 70
rect 369 53 371 58
rect 365 52 371 53
rect 369 47 371 52
rect 368 33 371 47
rect 294 18 300 21
rect 314 18 320 21
rect 334 18 340 29
rect 369 29 371 33
rect 374 42 380 53
rect 379 36 380 42
rect 374 33 380 36
rect 383 33 387 53
rect 404 50 408 53
rect 404 33 408 45
rect 384 29 385 33
rect 393 29 394 33
rect 354 25 358 27
rect 354 21 355 25
rect 393 18 397 29
rect 411 25 415 67
rect 464 59 470 70
rect 429 53 430 58
rect 427 50 430 53
rect 427 33 430 45
rect 449 53 450 58
rect 435 40 439 53
rect 438 35 439 40
rect 435 33 439 35
rect 445 33 450 53
rect 453 53 455 59
rect 479 54 480 59
rect 453 39 457 53
rect 453 33 458 34
rect 476 33 480 48
rect 453 29 455 33
rect 479 29 480 33
rect 405 21 414 25
rect 464 18 470 29
rect 247 11 334 18
rect 350 14 364 18
rect 368 14 388 18
rect 350 11 388 14
rect 400 14 424 18
rect 428 14 434 18
rect 400 12 434 14
rect 442 12 487 18
rect 400 11 487 12
rect 247 10 487 11
<< m2contact >>
rect 346 48 351 53
rect 364 47 369 52
rect 353 27 358 32
rect 374 36 379 42
rect 403 45 408 50
rect 425 45 430 50
rect 433 35 438 40
rect 453 34 458 39
rect 464 36 469 41
<< pm12contact >>
rect 370 62 375 67
rect 380 62 385 67
rect 300 36 305 46
rect 309 36 314 46
rect 338 39 343 44
rect 360 36 365 41
rect 390 36 395 41
rect 370 21 375 26
rect 380 21 385 26
rect 400 21 405 26
rect 430 62 435 67
rect 440 62 445 67
rect 419 36 424 41
rect 460 45 465 50
rect 430 21 435 26
rect 439 21 444 26
<< pdm12contact >>
rect 304 50 310 67
rect 324 59 330 67
rect 444 53 449 58
<< ndm12contact >>
rect 304 21 310 32
rect 324 21 330 27
<< metal2 >>
rect 371 72 446 75
rect 371 71 440 72
rect 371 67 376 71
rect 375 62 376 67
rect 390 62 430 67
rect 435 62 436 67
rect 371 59 376 62
rect 324 46 330 59
rect 351 48 364 52
rect 347 47 364 48
rect 373 51 376 59
rect 432 58 436 62
rect 450 58 456 62
rect 432 54 440 58
rect 373 47 386 51
rect 305 36 309 46
rect 314 36 330 46
rect 284 18 290 31
rect 324 27 330 36
rect 338 32 343 39
rect 365 36 374 41
rect 338 27 353 32
rect 383 26 386 47
rect 408 45 425 50
rect 434 49 440 54
rect 449 53 456 58
rect 434 44 448 49
rect 395 36 405 39
rect 391 35 405 36
rect 424 36 433 40
rect 419 35 433 36
rect 443 39 448 44
rect 385 21 386 26
rect 400 26 405 35
rect 443 34 453 39
rect 458 36 464 39
rect 458 34 469 36
rect 443 26 448 34
rect 444 21 448 26
rect 284 17 291 18
rect 284 11 310 17
rect 304 8 310 11
<< m3contact >>
rect 440 67 445 72
rect 294 50 304 67
rect 385 62 390 67
rect 294 21 304 32
rect 365 21 370 26
rect 425 21 430 26
<< m123contact >>
rect 450 62 456 67
rect 474 48 480 54
<< metal3 >>
rect 450 67 456 77
rect 259 42 265 59
rect 285 47 294 67
rect 380 62 385 67
rect 381 51 385 62
rect 440 54 446 67
rect 269 38 294 47
rect 275 36 294 38
rect 285 21 294 36
rect 371 46 385 51
rect 425 48 474 54
rect 371 26 376 46
rect 370 21 376 26
rect 425 26 431 48
rect 285 16 304 21
rect 285 14 484 16
rect 247 8 255 14
rect 285 10 487 14
rect 478 8 487 10
<< m345contact >>
rect 259 59 266 66
<< metal5 >>
rect 247 59 259 66
rect 266 59 487 66
use and  and_0
timestamp 1575783955
transform 1 0 251 0 1 6
box 0 4 42 72
<< labels >>
rlabel metal1 485 74 485 74 7 Vdd
rlabel metal5 253 62 253 62 1 y
rlabel metal2 307 9 307 9 1 z
rlabel pm12contact 463 47 463 47 1 clk
rlabel metal1 448 43 448 43 1 D
rlabel metal1 377 12 377 12 1 Gnd
rlabel metal1 365 74 365 74 1 Vdd
rlabel polycontact 323 42 323 42 1 Q
<< end >>
