magic
tech scmos
timestamp 1576184507
<< metal6 >>
rect 4063 19787 4297 20241
rect 5004 19805 5238 20259
rect 5890 19777 6124 20231
rect 6785 19796 7019 20250
rect 7693 19773 7927 20227
rect 8551 19782 8785 20236
rect 9460 19787 9694 20241
rect 10350 19805 10584 20259
rect 11236 19796 11470 20250
rect 12117 19796 12351 20250
rect 12998 19777 13232 20231
rect 13907 19764 14141 20218
rect 14747 19782 14981 20236
rect 16559 20126 20562 20373
rect 16559 19632 16806 20126
rect 20315 16434 20562 20126
rect 19509 16158 20562 16434
rect 20315 16152 20562 16158
rect -381 14386 97 14509
rect 19632 14394 19993 14457
rect -368 13526 110 13649
rect 19639 13531 19993 13594
rect -336 12634 142 12757
rect 19627 12649 19995 12712
rect -186 11748 112 11811
rect 19636 11740 19996 11803
rect 19634 10863 19999 10926
rect 19627 9997 20002 10060
rect 19636 9079 20005 9142
rect 19625 8199 20008 8262
rect 19641 6462 20016 6525
rect 19632 5549 20017 5612
rect 19627 4655 19922 4718
rect -1715 3938 -304 3948
rect -1715 3738 216 3938
rect -1715 3718 -304 3738
rect -1715 -815 -1485 3718
rect 4129 -815 4359 226
rect 5083 -179 5138 69
rect 5971 -184 6026 64
rect 6891 -175 6946 73
rect 7786 -200 7841 48
rect 8647 -192 8702 56
rect 9534 -208 9589 40
rect 10396 -208 10451 40
rect 11315 -208 11370 40
rect 12171 -419 12234 73
rect 12963 -75 13026 55
rect 13899 -52 13962 55
rect 12963 -138 13030 -75
rect 13760 -100 13962 -52
rect 14963 -71 15026 41
rect 14963 -92 15040 -71
rect 13760 -115 14520 -100
rect 13760 -138 13823 -115
rect 12967 -304 13030 -138
rect 13895 -163 14520 -115
rect 14975 -138 15040 -92
rect 12967 -367 13411 -304
rect 13348 -427 13411 -367
rect 14457 -437 14520 -163
rect 14977 -234 15040 -138
rect 14977 -297 15748 -234
rect 15685 -427 15748 -297
rect -1715 -1045 4359 -815
use ninepf  ninepf_16
timestamp 1085807705
transform -1 0 -238 0 -1 12245
box -52 60 3722 857
use chip  chip_0
timestamp 1576183136
transform 1 0 3013 0 1 17237
box -3013 -17237 16677 2672
use ninepf  ninepf_11
timestamp 1085807705
transform 1 0 20045 0 1 13965
box -52 60 3722 857
use ninepf  ninepf_10
timestamp 1085807705
transform 1 0 20045 0 1 13097
box -52 60 3722 857
use ninepf  ninepf_9
timestamp 1085807705
transform 1 0 20047 0 1 12220
box -52 60 3722 857
use ninepf  ninepf_8
timestamp 1085807705
transform 1 0 20048 0 1 11311
box -52 60 3722 857
use ninepf  ninepf_7
timestamp 1085807705
transform 1 0 20051 0 1 10434
box -52 60 3722 857
use ninepf  ninepf_6
timestamp 1085807705
transform 1 0 20054 0 1 9563
box -52 60 3722 857
use ninepf  ninepf_5
timestamp 1085807705
transform 1 0 20057 0 1 8650
box -52 60 3722 857
use ninepf  ninepf_4
timestamp 1085807705
transform 1 0 20060 0 1 7770
box -52 60 3722 857
use ninepf  ninepf_2
timestamp 1085807705
transform 1 0 20068 0 1 6031
box -52 60 3722 857
use ninepf  ninepf_1
timestamp 1085807705
transform 1 0 20069 0 1 5115
box -52 60 3722 857
use ninepf  ninepf_0
timestamp 1085807705
transform 1 0 19974 0 1 4226
box -52 60 3722 857
use ninepf  ninepf_12
timestamp 1085807705
transform 0 1 11737 -1 0 -471
box -52 60 3722 857
use ninepf  ninepf_13
timestamp 1085807705
transform 0 1 12914 -1 0 -479
box -52 60 3722 857
use ninepf  ninepf_14
timestamp 1085807705
transform 0 1 14028 -1 0 -489
box -52 60 3722 857
use ninepf  ninepf_15
timestamp 1085807705
transform 0 1 15251 -1 0 -479
box -52 60 3722 857
<< labels >>
rlabel metal6 12207 -230 12207 -230 1 c1
rlabel metal6 13136 -356 13136 -356 1 c2
rlabel metal6 14490 -331 14490 -331 1 c3
rlabel metal6 15716 -357 15716 -357 1 c4
rlabel metal6 19784 4686 19784 4686 1 c5
rlabel metal6 19828 5577 19828 5577 1 c6
rlabel metal6 19828 6494 19828 6494 1 c7
rlabel metal6 -107 11784 -107 11784 1 c0
rlabel metal6 19830 8226 19830 8226 1 d7
rlabel metal6 19816 9108 19816 9108 1 d6
rlabel metal6 19848 10023 19848 10023 1 d5
rlabel metal6 19816 10899 19816 10899 1 d4
rlabel metal6 19781 11768 19781 11768 1 d3
rlabel metal6 19799 12681 19799 12681 1 d2
rlabel metal6 19789 13563 19789 13563 1 d1
rlabel metal6 19785 14425 19785 14425 1 d0
rlabel metal6 5109 -104 5109 -104 1 opcode0
rlabel metal6 6009 -96 6009 -96 1 cen
rlabel metal6 6919 -79 6919 -79 1 opcode1
rlabel metal6 7813 -100 7813 -100 1 den
rlabel metal6 8671 -94 8671 -94 1 b5
rlabel metal6 9563 -106 9563 -106 1 opcode2
rlabel metal6 10423 -106 10423 -106 1 b6
rlabel metal6 11348 -127 11348 -127 1 b7
rlabel metal6 -239 12694 -239 12694 1 clk
rlabel metal6 -262 13582 -262 13582 1 bctrl
rlabel metal6 -264 14450 -264 14450 1 actrl
rlabel metal6 4172 20069 4172 20069 1 b4
rlabel metal6 5147 20069 5147 20069 1 b3
rlabel metal6 6021 20085 6021 20085 1 b2
rlabel metal6 6918 20057 6918 20057 1 b1
rlabel metal6 7813 20048 7813 20048 1 b0
rlabel metal6 8659 20036 8659 20036 1 a0
rlabel metal6 9589 20045 9589 20045 1 a1
rlabel metal6 10468 20043 10468 20043 1 a2
rlabel metal6 11349 20027 11349 20027 1 a3
rlabel metal6 12234 20038 12234 20038 1 a4
rlabel metal6 13106 20052 13106 20052 1 a5
rlabel metal6 14026 20036 14026 20036 1 a6
rlabel metal6 14861 20043 14861 20043 1 a7
rlabel metal6 20404 16300 20404 16300 1 Vdd
rlabel metal6 -624 3818 -624 3828 1 Gnd
<< end >>
