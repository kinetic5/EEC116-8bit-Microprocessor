magic
tech scmos
timestamp 1575998097
<< metal1 >>
rect -1773 1214 15766 1543
rect -1773 -15993 -1444 1214
rect -1216 657 15202 986
rect -1216 -15423 -887 657
rect 232 650 561 657
rect 232 456 561 457
rect -667 127 14661 456
rect -666 -14873 -337 127
rect -116 -95 213 -94
rect 577 -95 14100 -94
rect -116 -423 14100 -95
rect -116 -14336 213 -423
rect 13771 -3679 14100 -423
rect 13756 -4525 14100 -3679
rect 13756 -14336 14085 -4525
rect -116 -14341 222 -14336
rect 582 -14341 14085 -14336
rect -116 -14658 14085 -14341
rect -116 -14665 222 -14658
rect 588 -14665 14085 -14658
rect 14323 -14871 14655 127
rect 14873 -1424 15202 657
rect 232 -14873 561 -14872
rect 866 -14873 14655 -14871
rect -666 -15200 14655 -14873
rect 14870 -3055 15202 -1424
rect -666 -15202 14649 -15200
rect -664 -15211 14649 -15202
rect 232 -15423 561 -15420
rect 14870 -15423 15199 -3055
rect 15437 -14766 15766 1214
rect -1216 -15752 15199 -15423
rect 15521 -14769 15766 -14766
rect 15521 -15983 15646 -14769
rect 15437 -15989 15646 -15983
rect 15437 -15993 15768 -15989
rect -1773 -15998 8414 -15993
rect -1773 -16081 14470 -15998
rect -1773 -16210 15766 -16081
rect -1773 -16322 14469 -16210
rect 7835 -16324 14469 -16322
rect 15753 -16324 15766 -16210
rect 7835 -16327 15766 -16324
<< metal2 >>
rect 240 1543 15763 1546
rect -1774 1217 15763 1543
rect -1774 1214 890 1217
rect -1774 -15992 -1445 1214
rect -929 981 15213 982
rect -1217 653 15213 981
rect -1217 652 896 653
rect -1217 -15428 -888 652
rect -667 444 876 457
rect -667 129 14649 444
rect -667 -14883 -339 129
rect 467 116 14649 129
rect 1720 -95 2049 -94
rect 2520 -95 14096 -93
rect -116 -422 14096 -95
rect -116 -423 3442 -422
rect -116 -424 222 -423
rect 582 -424 3442 -423
rect -116 -14333 213 -424
rect 13767 -14333 14096 -422
rect -116 -14341 222 -14333
rect 582 -14341 14096 -14333
rect -116 -14662 14096 -14341
rect 14321 -14883 14649 116
rect -667 -15211 14649 -14883
rect 14884 -15428 15213 653
rect -1217 -15757 15213 -15428
rect 15434 -14766 15763 1217
rect 15521 -14769 15763 -14766
rect 15521 -14771 15646 -14769
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -15986 15646 -14771
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -15993 15768 -15992
rect -1774 -16081 14470 -15993
rect -1774 -16090 15763 -16081
rect -1774 -16204 14468 -16090
rect 15752 -16204 15763 -16090
rect -1774 -16210 15763 -16204
rect -1774 -16321 14469 -16210
rect 15753 -16321 15763 -16210
<< m123contact >>
rect 15434 -15983 15521 -14766
rect 15646 -15989 15768 -14799
rect 14470 -16081 15768 -15993
rect 14469 -16324 15753 -16210
<< metal3 >>
rect -1774 1217 15763 1546
rect -1774 -15992 -1445 1217
rect -1224 982 1544 984
rect -1224 655 15213 982
rect -1224 -15428 -895 655
rect 466 653 15213 655
rect -667 444 1547 454
rect -667 125 14656 444
rect -667 -14889 -338 125
rect 108 115 14656 125
rect -115 -101 2593 -94
rect -115 -423 14094 -101
rect -115 -14334 214 -423
rect 2416 -430 14094 -423
rect 13765 -14334 14094 -430
rect -115 -14663 14094 -14334
rect 14327 -14889 14656 115
rect -667 -15218 14656 -14889
rect 14884 -15428 15213 653
rect -1224 -15757 15213 -15428
rect 15434 -14766 15763 1217
rect 15521 -14769 15763 -14766
rect 15521 -14771 15646 -14769
rect 15521 -15983 15529 -14771
rect 15434 -15986 15529 -15983
rect 15644 -15986 15646 -14771
rect 15434 -15989 15646 -15986
rect 15434 -15992 15768 -15989
rect -1774 -15993 15768 -15992
rect -1774 -16081 14470 -15993
rect -1774 -16090 15763 -16081
rect -1774 -16204 14468 -16090
rect 15752 -16204 15763 -16090
rect -1774 -16210 15763 -16204
rect -1774 -16321 14469 -16210
rect 15753 -16321 15763 -16210
<< m234contact >>
rect 15529 -15986 15644 -14771
rect 14468 -16204 15752 -16090
<< metal4 >>
rect 1879 1539 15433 1549
rect 15529 1539 15770 1549
rect -1767 1220 15770 1539
rect -1767 1210 8012 1220
rect -1767 -15992 -1438 1210
rect -1217 984 2672 989
rect -1217 660 15213 984
rect -1217 -15415 -888 660
rect 1910 655 15213 660
rect -667 451 2201 454
rect -667 125 14656 451
rect -667 -14882 -338 125
rect -322 122 14656 125
rect -115 -94 6919 -87
rect -115 -416 14094 -94
rect -115 -14334 214 -416
rect 2735 -423 14094 -416
rect 13765 -14334 14094 -423
rect -115 -14663 14094 -14334
rect 14327 -14882 14656 122
rect -667 -15211 14656 -14882
rect 14884 -15415 15213 655
rect -1217 -15744 15213 -15415
rect 15433 -14771 15762 1220
rect 15433 -15986 15529 -14771
rect 15644 -15986 15762 -14771
rect 15433 -15989 15762 -15986
rect 15433 -15992 15768 -15989
rect -1788 -15993 15768 -15992
rect -1788 -16090 15762 -15993
rect -1788 -16204 14468 -16090
rect 15752 -16204 15762 -16090
rect -1788 -16321 15762 -16204
use pad  pad_48
timestamp 1575998002
transform 1 0 -29 0 1 2000
box -3 -4 672 668
use pad  pad_49
timestamp 1575998002
transform 1 0 860 0 1 2000
box -3 -4 672 668
use pad  pad_50
timestamp 1575998002
transform 1 0 1749 0 1 2000
box -3 -4 672 668
use pad  pad_51
timestamp 1575998002
transform 1 0 2638 0 1 2000
box -3 -4 672 668
use pad  pad_52
timestamp 1575998002
transform 1 0 3527 0 1 2000
box -3 -4 672 668
use pad  pad_53
timestamp 1575998002
transform 1 0 4416 0 1 2000
box -3 -4 672 668
use pad  pad_54
timestamp 1575998002
transform 1 0 5305 0 1 2000
box -3 -4 672 668
use pad  pad_55
timestamp 1575998002
transform 1 0 6194 0 1 2000
box -3 -4 672 668
use pad  pad_56
timestamp 1575998002
transform 1 0 7083 0 1 2000
box -3 -4 672 668
use pad  pad_57
timestamp 1575998002
transform 1 0 7972 0 1 2000
box -3 -4 672 668
use pad  pad_58
timestamp 1575998002
transform 1 0 8861 0 1 2000
box -3 -4 672 668
use pad  pad_59
timestamp 1575998002
transform 1 0 9750 0 1 2000
box -3 -4 672 668
use pad  pad_60
timestamp 1575998002
transform 1 0 10639 0 1 2000
box -3 -4 672 668
use pad  pad_61
timestamp 1575998002
transform 1 0 11528 0 1 2000
box -3 -4 672 668
use pad  pad_62
timestamp 1575998002
transform 1 0 12417 0 1 2000
box -3 -4 672 668
use pad  pad_63
timestamp 1575998002
transform 1 0 13306 0 1 2000
box -3 -4 672 668
use pad  pad_32
timestamp 1575998002
transform 0 1 -2998 -1 0 -662
box -3 -4 672 668
use pad  pad_16
timestamp 1575998002
transform 0 1 16001 -1 0 -645
box -3 -4 672 668
use pad  pad_33
timestamp 1575998002
transform 0 1 -2998 -1 0 -1551
box -3 -4 672 668
use pad  pad_17
timestamp 1575998002
transform 0 1 16001 -1 0 -1534
box -3 -4 672 668
use pad  pad_34
timestamp 1575998002
transform 0 1 -2998 -1 0 -2440
box -3 -4 672 668
use pad  pad_18
timestamp 1575998002
transform 0 1 16001 -1 0 -2423
box -3 -4 672 668
use pad  pad_35
timestamp 1575998002
transform 0 1 -2998 -1 0 -3329
box -3 -4 672 668
use pad  pad_19
timestamp 1575998002
transform 0 1 16001 -1 0 -3312
box -3 -4 672 668
use pad  pad_36
timestamp 1575998002
transform 0 1 -2998 -1 0 -4218
box -3 -4 672 668
use pad  pad_20
timestamp 1575998002
transform 0 1 16001 -1 0 -4201
box -3 -4 672 668
use pad  pad_37
timestamp 1575998002
transform 0 1 -2998 -1 0 -5107
box -3 -4 672 668
use pad  pad_21
timestamp 1575998002
transform 0 1 16001 -1 0 -5090
box -3 -4 672 668
use pad  pad_38
timestamp 1575998002
transform 0 1 -2998 -1 0 -5996
box -3 -4 672 668
use pad  pad_22
timestamp 1575998002
transform 0 1 16001 -1 0 -5979
box -3 -4 672 668
use pad  pad_39
timestamp 1575998002
transform 0 1 -2998 -1 0 -6885
box -3 -4 672 668
use pad  pad_23
timestamp 1575998002
transform 0 1 16001 -1 0 -6868
box -3 -4 672 668
use pad  pad_40
timestamp 1575998002
transform 0 1 -2998 -1 0 -7774
box -3 -4 672 668
use pad  pad_24
timestamp 1575998002
transform 0 1 16001 -1 0 -7757
box -3 -4 672 668
use pad  pad_41
timestamp 1575998002
transform 0 1 -2998 -1 0 -8663
box -3 -4 672 668
use pad  pad_25
timestamp 1575998002
transform 0 1 16001 -1 0 -8646
box -3 -4 672 668
use pad  pad_42
timestamp 1575998002
transform 0 1 -2998 -1 0 -9552
box -3 -4 672 668
use pad  pad_26
timestamp 1575998002
transform 0 1 16001 -1 0 -9535
box -3 -4 672 668
use pad  pad_43
timestamp 1575998002
transform 0 1 -2998 -1 0 -10441
box -3 -4 672 668
use pad  pad_27
timestamp 1575998002
transform 0 1 16001 -1 0 -10424
box -3 -4 672 668
use pad  pad_44
timestamp 1575998002
transform 0 1 -2998 -1 0 -11330
box -3 -4 672 668
use pad  pad_28
timestamp 1575998002
transform 0 1 16001 -1 0 -11313
box -3 -4 672 668
use pad  pad_45
timestamp 1575998002
transform 0 1 -2998 -1 0 -12219
box -3 -4 672 668
use pad  pad_29
timestamp 1575998002
transform 0 1 16001 -1 0 -12202
box -3 -4 672 668
use pad  pad_46
timestamp 1575998002
transform 0 1 -2998 -1 0 -13108
box -3 -4 672 668
use pad  pad_30
timestamp 1575998002
transform 0 1 16001 -1 0 -13091
box -3 -4 672 668
use pad  pad_47
timestamp 1575998002
transform 0 1 -2998 -1 0 -13997
box -3 -4 672 668
use pad  pad_31
timestamp 1575998002
transform 0 1 16001 -1 0 -13980
box -3 -4 672 668
use pad  pad_0
timestamp 1575998002
transform 1 0 0 0 1 -17223
box -3 -4 672 668
use pad  pad_1
timestamp 1575998002
transform 1 0 889 0 1 -17223
box -3 -4 672 668
use pad  pad_2
timestamp 1575998002
transform 1 0 1778 0 1 -17223
box -3 -4 672 668
use pad  pad_3
timestamp 1575998002
transform 1 0 2667 0 1 -17223
box -3 -4 672 668
use pad  pad_4
timestamp 1575998002
transform 1 0 3556 0 1 -17223
box -3 -4 672 668
use pad  pad_5
timestamp 1575998002
transform 1 0 4445 0 1 -17223
box -3 -4 672 668
use pad  pad_6
timestamp 1575998002
transform 1 0 5334 0 1 -17223
box -3 -4 672 668
use pad  pad_7
timestamp 1575998002
transform 1 0 6223 0 1 -17223
box -3 -4 672 668
use pad  pad_8
timestamp 1575998002
transform 1 0 7112 0 1 -17223
box -3 -4 672 668
use pad  pad_9
timestamp 1575998002
transform 1 0 8001 0 1 -17223
box -3 -4 672 668
use pad  pad_10
timestamp 1575998002
transform 1 0 8890 0 1 -17223
box -3 -4 672 668
use pad  pad_11
timestamp 1575998002
transform 1 0 9779 0 1 -17223
box -3 -4 672 668
use pad  pad_12
timestamp 1575998002
transform 1 0 10668 0 1 -17223
box -3 -4 672 668
use pad  pad_13
timestamp 1575998002
transform 1 0 11557 0 1 -17223
box -3 -4 672 668
use pad  pad_14
timestamp 1575998002
transform 1 0 12446 0 1 -17223
box -3 -4 672 668
use pad  pad_15
timestamp 1575998002
transform 1 0 13335 0 1 -17223
box -3 -4 672 668
<< labels >>
rlabel metal4 6989 -16182 6989 -16182 1 VddIo
rlabel metal4 7131 -15637 7131 -15637 1 GndIo
rlabel metal4 7143 -15058 7143 -15058 1 VddCore
rlabel metal4 7143 -14490 7143 -14490 1 GndCore
<< end >>
