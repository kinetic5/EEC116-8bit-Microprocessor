magic
tech scmos
timestamp 1575762367
<< ntransistor >>
rect -7 -141 -5 -137
rect 3 -141 5 -137
<< ptransistor >>
rect -7 -117 -5 -111
rect 3 -117 5 -111
<< ndiffusion >>
rect -8 -141 -7 -137
rect -5 -141 -4 -137
rect 2 -141 3 -137
rect 5 -141 6 -137
<< pdiffusion >>
rect -8 -117 -7 -111
rect -5 -117 -3 -111
rect 1 -117 3 -111
rect 5 -112 10 -111
rect 5 -117 6 -112
<< ndcontact >>
rect -12 -141 -8 -137
rect -4 -141 2 -137
rect 6 -141 10 -137
<< pdcontact >>
rect -12 -117 -8 -111
rect -3 -117 1 -111
rect 6 -117 10 -112
<< polysilicon >>
rect -7 -111 -5 -108
rect 3 -111 5 -108
rect -7 -124 -5 -117
rect 3 -124 5 -117
rect -7 -137 -5 -130
rect 3 -137 5 -130
rect -7 -144 -5 -141
rect 3 -144 5 -141
<< metal1 >>
rect -13 -100 13 -92
rect 130 -97 132 -95
rect -13 -117 -12 -111
rect -13 -137 -10 -117
rect -3 -132 1 -117
rect 5 -117 6 -112
rect 5 -132 8 -117
rect 180 -125 183 -121
rect -13 -141 -12 -137
rect 5 -141 6 -132
rect -13 -160 13 -152
rect 118 -159 120 -157
<< m2contact >>
rect -3 -137 2 -132
rect 6 -137 11 -132
<< pm12contact >>
rect -9 -108 -4 -103
rect 1 -108 6 -103
rect -9 -149 -4 -144
rect 1 -149 6 -144
<< metal2 >>
rect 30 -92 35 -89
rect 1 -116 6 -108
rect -2 -117 6 -116
rect -11 -119 6 -117
rect 41 -117 49 -112
rect -11 -120 1 -119
rect -11 -129 -7 -120
rect -10 -144 -7 -129
rect -3 -128 5 -125
rect 41 -126 44 -117
rect -3 -132 2 -128
rect -10 -149 -9 -144
rect 11 -153 16 -132
rect 179 -153 184 -129
rect 11 -157 184 -153
<< m3contact >>
rect -11 -113 -6 -108
rect 5 -128 10 -123
rect 40 -131 45 -126
rect 1 -154 6 -149
<< metal3 >>
rect -9 -108 -4 -103
rect -6 -113 -4 -108
rect -9 -144 -4 -113
rect 10 -128 40 -126
rect 5 -131 40 -128
rect -9 -149 6 -144
use DFF  DFF_0
timestamp 1575762319
transform 1 0 119 0 1 -128
box -108 -32 68 36
<< labels >>
rlabel metal1 -12 -132 -12 -132 1 D
rlabel pm12contact -6 -146 -6 -146 1 EN
rlabel metal3 3 -146 3 -146 1 ENbar
rlabel metal2 32 -91 32 -91 5 clk
rlabel metal2 182 -132 182 -132 7 Q
rlabel metal1 182 -123 182 -123 7 Qbar
rlabel metal1 119 -158 119 -158 1 Gnd
rlabel metal1 131 -96 131 -96 1 Vdd
<< end >>
